module compressorInput(
  output [11:0] io_input_currentByteOut,
  input  [7:0]  io_input_dataIn_0,
  input         io_input_valid,
  output        io_input_ready,
  input  [11:0] io_currentByte,
  input         io_dataOut_ready,
  output        io_dataOut_valid,
  output [7:0]  io_dataOut_bits_0
);
  assign io_input_currentByteOut = io_currentByte; // @[compressorInput.scala 63:29]
  assign io_input_ready = io_dataOut_ready; // @[compressorInput.scala 31:20]
  assign io_dataOut_valid = io_input_valid; // @[compressorInput.scala 61:22]
  assign io_dataOut_bits_0 = io_input_dataIn_0; // @[compressorInput.scala 62:21]
endmodule
module characterFrequencyCounter(
  input         clock,
  input         reset,
  input         io_start,
  output        io_dataIn_ready,
  input  [7:0]  io_dataIn_bits_0,
  output [11:0] io_currentByte,
  output [12:0] io_frequencies_0,
  output [12:0] io_frequencies_1,
  output [12:0] io_frequencies_2,
  output [12:0] io_frequencies_3,
  output [12:0] io_frequencies_4,
  output [12:0] io_frequencies_5,
  output [12:0] io_frequencies_6,
  output [12:0] io_frequencies_7,
  output [12:0] io_frequencies_8,
  output [12:0] io_frequencies_9,
  output [12:0] io_frequencies_10,
  output [12:0] io_frequencies_11,
  output [12:0] io_frequencies_12,
  output [12:0] io_frequencies_13,
  output [12:0] io_frequencies_14,
  output [12:0] io_frequencies_15,
  output [12:0] io_frequencies_16,
  output [12:0] io_frequencies_17,
  output [12:0] io_frequencies_18,
  output [12:0] io_frequencies_19,
  output [12:0] io_frequencies_20,
  output [12:0] io_frequencies_21,
  output [12:0] io_frequencies_22,
  output [12:0] io_frequencies_23,
  output [12:0] io_frequencies_24,
  output [12:0] io_frequencies_25,
  output [12:0] io_frequencies_26,
  output [12:0] io_frequencies_27,
  output [12:0] io_frequencies_28,
  output [12:0] io_frequencies_29,
  output [12:0] io_frequencies_30,
  output [12:0] io_frequencies_31,
  output [12:0] io_frequencies_32,
  output [12:0] io_frequencies_33,
  output [12:0] io_frequencies_34,
  output [12:0] io_frequencies_35,
  output [12:0] io_frequencies_36,
  output [12:0] io_frequencies_37,
  output [12:0] io_frequencies_38,
  output [12:0] io_frequencies_39,
  output [12:0] io_frequencies_40,
  output [12:0] io_frequencies_41,
  output [12:0] io_frequencies_42,
  output [12:0] io_frequencies_43,
  output [12:0] io_frequencies_44,
  output [12:0] io_frequencies_45,
  output [12:0] io_frequencies_46,
  output [12:0] io_frequencies_47,
  output [12:0] io_frequencies_48,
  output [12:0] io_frequencies_49,
  output [12:0] io_frequencies_50,
  output [12:0] io_frequencies_51,
  output [12:0] io_frequencies_52,
  output [12:0] io_frequencies_53,
  output [12:0] io_frequencies_54,
  output [12:0] io_frequencies_55,
  output [12:0] io_frequencies_56,
  output [12:0] io_frequencies_57,
  output [12:0] io_frequencies_58,
  output [12:0] io_frequencies_59,
  output [12:0] io_frequencies_60,
  output [12:0] io_frequencies_61,
  output [12:0] io_frequencies_62,
  output [12:0] io_frequencies_63,
  output [12:0] io_frequencies_64,
  output [12:0] io_frequencies_65,
  output [12:0] io_frequencies_66,
  output [12:0] io_frequencies_67,
  output [12:0] io_frequencies_68,
  output [12:0] io_frequencies_69,
  output [12:0] io_frequencies_70,
  output [12:0] io_frequencies_71,
  output [12:0] io_frequencies_72,
  output [12:0] io_frequencies_73,
  output [12:0] io_frequencies_74,
  output [12:0] io_frequencies_75,
  output [12:0] io_frequencies_76,
  output [12:0] io_frequencies_77,
  output [12:0] io_frequencies_78,
  output [12:0] io_frequencies_79,
  output [12:0] io_frequencies_80,
  output [12:0] io_frequencies_81,
  output [12:0] io_frequencies_82,
  output [12:0] io_frequencies_83,
  output [12:0] io_frequencies_84,
  output [12:0] io_frequencies_85,
  output [12:0] io_frequencies_86,
  output [12:0] io_frequencies_87,
  output [12:0] io_frequencies_88,
  output [12:0] io_frequencies_89,
  output [12:0] io_frequencies_90,
  output [12:0] io_frequencies_91,
  output [12:0] io_frequencies_92,
  output [12:0] io_frequencies_93,
  output [12:0] io_frequencies_94,
  output [12:0] io_frequencies_95,
  output [12:0] io_frequencies_96,
  output [12:0] io_frequencies_97,
  output [12:0] io_frequencies_98,
  output [12:0] io_frequencies_99,
  output [12:0] io_frequencies_100,
  output [12:0] io_frequencies_101,
  output [12:0] io_frequencies_102,
  output [12:0] io_frequencies_103,
  output [12:0] io_frequencies_104,
  output [12:0] io_frequencies_105,
  output [12:0] io_frequencies_106,
  output [12:0] io_frequencies_107,
  output [12:0] io_frequencies_108,
  output [12:0] io_frequencies_109,
  output [12:0] io_frequencies_110,
  output [12:0] io_frequencies_111,
  output [12:0] io_frequencies_112,
  output [12:0] io_frequencies_113,
  output [12:0] io_frequencies_114,
  output [12:0] io_frequencies_115,
  output [12:0] io_frequencies_116,
  output [12:0] io_frequencies_117,
  output [12:0] io_frequencies_118,
  output [12:0] io_frequencies_119,
  output [12:0] io_frequencies_120,
  output [12:0] io_frequencies_121,
  output [12:0] io_frequencies_122,
  output [12:0] io_frequencies_123,
  output [12:0] io_frequencies_124,
  output [12:0] io_frequencies_125,
  output [12:0] io_frequencies_126,
  output [12:0] io_frequencies_127,
  output [12:0] io_frequencies_128,
  output [12:0] io_frequencies_129,
  output [12:0] io_frequencies_130,
  output [12:0] io_frequencies_131,
  output [12:0] io_frequencies_132,
  output [12:0] io_frequencies_133,
  output [12:0] io_frequencies_134,
  output [12:0] io_frequencies_135,
  output [12:0] io_frequencies_136,
  output [12:0] io_frequencies_137,
  output [12:0] io_frequencies_138,
  output [12:0] io_frequencies_139,
  output [12:0] io_frequencies_140,
  output [12:0] io_frequencies_141,
  output [12:0] io_frequencies_142,
  output [12:0] io_frequencies_143,
  output [12:0] io_frequencies_144,
  output [12:0] io_frequencies_145,
  output [12:0] io_frequencies_146,
  output [12:0] io_frequencies_147,
  output [12:0] io_frequencies_148,
  output [12:0] io_frequencies_149,
  output [12:0] io_frequencies_150,
  output [12:0] io_frequencies_151,
  output [12:0] io_frequencies_152,
  output [12:0] io_frequencies_153,
  output [12:0] io_frequencies_154,
  output [12:0] io_frequencies_155,
  output [12:0] io_frequencies_156,
  output [12:0] io_frequencies_157,
  output [12:0] io_frequencies_158,
  output [12:0] io_frequencies_159,
  output [12:0] io_frequencies_160,
  output [12:0] io_frequencies_161,
  output [12:0] io_frequencies_162,
  output [12:0] io_frequencies_163,
  output [12:0] io_frequencies_164,
  output [12:0] io_frequencies_165,
  output [12:0] io_frequencies_166,
  output [12:0] io_frequencies_167,
  output [12:0] io_frequencies_168,
  output [12:0] io_frequencies_169,
  output [12:0] io_frequencies_170,
  output [12:0] io_frequencies_171,
  output [12:0] io_frequencies_172,
  output [12:0] io_frequencies_173,
  output [12:0] io_frequencies_174,
  output [12:0] io_frequencies_175,
  output [12:0] io_frequencies_176,
  output [12:0] io_frequencies_177,
  output [12:0] io_frequencies_178,
  output [12:0] io_frequencies_179,
  output [12:0] io_frequencies_180,
  output [12:0] io_frequencies_181,
  output [12:0] io_frequencies_182,
  output [12:0] io_frequencies_183,
  output [12:0] io_frequencies_184,
  output [12:0] io_frequencies_185,
  output [12:0] io_frequencies_186,
  output [12:0] io_frequencies_187,
  output [12:0] io_frequencies_188,
  output [12:0] io_frequencies_189,
  output [12:0] io_frequencies_190,
  output [12:0] io_frequencies_191,
  output [12:0] io_frequencies_192,
  output [12:0] io_frequencies_193,
  output [12:0] io_frequencies_194,
  output [12:0] io_frequencies_195,
  output [12:0] io_frequencies_196,
  output [12:0] io_frequencies_197,
  output [12:0] io_frequencies_198,
  output [12:0] io_frequencies_199,
  output [12:0] io_frequencies_200,
  output [12:0] io_frequencies_201,
  output [12:0] io_frequencies_202,
  output [12:0] io_frequencies_203,
  output [12:0] io_frequencies_204,
  output [12:0] io_frequencies_205,
  output [12:0] io_frequencies_206,
  output [12:0] io_frequencies_207,
  output [12:0] io_frequencies_208,
  output [12:0] io_frequencies_209,
  output [12:0] io_frequencies_210,
  output [12:0] io_frequencies_211,
  output [12:0] io_frequencies_212,
  output [12:0] io_frequencies_213,
  output [12:0] io_frequencies_214,
  output [12:0] io_frequencies_215,
  output [12:0] io_frequencies_216,
  output [12:0] io_frequencies_217,
  output [12:0] io_frequencies_218,
  output [12:0] io_frequencies_219,
  output [12:0] io_frequencies_220,
  output [12:0] io_frequencies_221,
  output [12:0] io_frequencies_222,
  output [12:0] io_frequencies_223,
  output [12:0] io_frequencies_224,
  output [12:0] io_frequencies_225,
  output [12:0] io_frequencies_226,
  output [12:0] io_frequencies_227,
  output [12:0] io_frequencies_228,
  output [12:0] io_frequencies_229,
  output [12:0] io_frequencies_230,
  output [12:0] io_frequencies_231,
  output [12:0] io_frequencies_232,
  output [12:0] io_frequencies_233,
  output [12:0] io_frequencies_234,
  output [12:0] io_frequencies_235,
  output [12:0] io_frequencies_236,
  output [12:0] io_frequencies_237,
  output [12:0] io_frequencies_238,
  output [12:0] io_frequencies_239,
  output [12:0] io_frequencies_240,
  output [12:0] io_frequencies_241,
  output [12:0] io_frequencies_242,
  output [12:0] io_frequencies_243,
  output [12:0] io_frequencies_244,
  output [12:0] io_frequencies_245,
  output [12:0] io_frequencies_246,
  output [12:0] io_frequencies_247,
  output [12:0] io_frequencies_248,
  output [12:0] io_frequencies_249,
  output [12:0] io_frequencies_250,
  output [12:0] io_frequencies_251,
  output [12:0] io_frequencies_252,
  output [12:0] io_frequencies_253,
  output [12:0] io_frequencies_254,
  output [12:0] io_frequencies_255,
  output        io_finished
);
  reg  state; // @[characterFrequencyCounter.scala 29:22]
  reg [31:0] _RAND_0;
  reg [12:0] currentByte; // @[characterFrequencyCounter.scala 33:24]
  reg [31:0] _RAND_1;
  reg [12:0] frequencyTotals_0; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_2;
  reg [12:0] frequencyTotals_1; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_3;
  reg [12:0] frequencyTotals_2; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_4;
  reg [12:0] frequencyTotals_3; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_5;
  reg [12:0] frequencyTotals_4; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_6;
  reg [12:0] frequencyTotals_5; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_7;
  reg [12:0] frequencyTotals_6; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_8;
  reg [12:0] frequencyTotals_7; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_9;
  reg [12:0] frequencyTotals_8; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_10;
  reg [12:0] frequencyTotals_9; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_11;
  reg [12:0] frequencyTotals_10; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_12;
  reg [12:0] frequencyTotals_11; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_13;
  reg [12:0] frequencyTotals_12; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_14;
  reg [12:0] frequencyTotals_13; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_15;
  reg [12:0] frequencyTotals_14; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_16;
  reg [12:0] frequencyTotals_15; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_17;
  reg [12:0] frequencyTotals_16; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_18;
  reg [12:0] frequencyTotals_17; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_19;
  reg [12:0] frequencyTotals_18; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_20;
  reg [12:0] frequencyTotals_19; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_21;
  reg [12:0] frequencyTotals_20; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_22;
  reg [12:0] frequencyTotals_21; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_23;
  reg [12:0] frequencyTotals_22; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_24;
  reg [12:0] frequencyTotals_23; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_25;
  reg [12:0] frequencyTotals_24; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_26;
  reg [12:0] frequencyTotals_25; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_27;
  reg [12:0] frequencyTotals_26; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_28;
  reg [12:0] frequencyTotals_27; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_29;
  reg [12:0] frequencyTotals_28; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_30;
  reg [12:0] frequencyTotals_29; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_31;
  reg [12:0] frequencyTotals_30; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_32;
  reg [12:0] frequencyTotals_31; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_33;
  reg [12:0] frequencyTotals_32; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_34;
  reg [12:0] frequencyTotals_33; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_35;
  reg [12:0] frequencyTotals_34; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_36;
  reg [12:0] frequencyTotals_35; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_37;
  reg [12:0] frequencyTotals_36; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_38;
  reg [12:0] frequencyTotals_37; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_39;
  reg [12:0] frequencyTotals_38; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_40;
  reg [12:0] frequencyTotals_39; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_41;
  reg [12:0] frequencyTotals_40; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_42;
  reg [12:0] frequencyTotals_41; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_43;
  reg [12:0] frequencyTotals_42; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_44;
  reg [12:0] frequencyTotals_43; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_45;
  reg [12:0] frequencyTotals_44; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_46;
  reg [12:0] frequencyTotals_45; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_47;
  reg [12:0] frequencyTotals_46; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_48;
  reg [12:0] frequencyTotals_47; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_49;
  reg [12:0] frequencyTotals_48; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_50;
  reg [12:0] frequencyTotals_49; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_51;
  reg [12:0] frequencyTotals_50; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_52;
  reg [12:0] frequencyTotals_51; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_53;
  reg [12:0] frequencyTotals_52; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_54;
  reg [12:0] frequencyTotals_53; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_55;
  reg [12:0] frequencyTotals_54; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_56;
  reg [12:0] frequencyTotals_55; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_57;
  reg [12:0] frequencyTotals_56; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_58;
  reg [12:0] frequencyTotals_57; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_59;
  reg [12:0] frequencyTotals_58; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_60;
  reg [12:0] frequencyTotals_59; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_61;
  reg [12:0] frequencyTotals_60; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_62;
  reg [12:0] frequencyTotals_61; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_63;
  reg [12:0] frequencyTotals_62; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_64;
  reg [12:0] frequencyTotals_63; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_65;
  reg [12:0] frequencyTotals_64; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_66;
  reg [12:0] frequencyTotals_65; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_67;
  reg [12:0] frequencyTotals_66; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_68;
  reg [12:0] frequencyTotals_67; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_69;
  reg [12:0] frequencyTotals_68; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_70;
  reg [12:0] frequencyTotals_69; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_71;
  reg [12:0] frequencyTotals_70; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_72;
  reg [12:0] frequencyTotals_71; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_73;
  reg [12:0] frequencyTotals_72; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_74;
  reg [12:0] frequencyTotals_73; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_75;
  reg [12:0] frequencyTotals_74; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_76;
  reg [12:0] frequencyTotals_75; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_77;
  reg [12:0] frequencyTotals_76; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_78;
  reg [12:0] frequencyTotals_77; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_79;
  reg [12:0] frequencyTotals_78; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_80;
  reg [12:0] frequencyTotals_79; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_81;
  reg [12:0] frequencyTotals_80; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_82;
  reg [12:0] frequencyTotals_81; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_83;
  reg [12:0] frequencyTotals_82; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_84;
  reg [12:0] frequencyTotals_83; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_85;
  reg [12:0] frequencyTotals_84; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_86;
  reg [12:0] frequencyTotals_85; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_87;
  reg [12:0] frequencyTotals_86; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_88;
  reg [12:0] frequencyTotals_87; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_89;
  reg [12:0] frequencyTotals_88; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_90;
  reg [12:0] frequencyTotals_89; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_91;
  reg [12:0] frequencyTotals_90; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_92;
  reg [12:0] frequencyTotals_91; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_93;
  reg [12:0] frequencyTotals_92; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_94;
  reg [12:0] frequencyTotals_93; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_95;
  reg [12:0] frequencyTotals_94; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_96;
  reg [12:0] frequencyTotals_95; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_97;
  reg [12:0] frequencyTotals_96; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_98;
  reg [12:0] frequencyTotals_97; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_99;
  reg [12:0] frequencyTotals_98; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_100;
  reg [12:0] frequencyTotals_99; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_101;
  reg [12:0] frequencyTotals_100; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_102;
  reg [12:0] frequencyTotals_101; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_103;
  reg [12:0] frequencyTotals_102; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_104;
  reg [12:0] frequencyTotals_103; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_105;
  reg [12:0] frequencyTotals_104; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_106;
  reg [12:0] frequencyTotals_105; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_107;
  reg [12:0] frequencyTotals_106; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_108;
  reg [12:0] frequencyTotals_107; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_109;
  reg [12:0] frequencyTotals_108; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_110;
  reg [12:0] frequencyTotals_109; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_111;
  reg [12:0] frequencyTotals_110; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_112;
  reg [12:0] frequencyTotals_111; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_113;
  reg [12:0] frequencyTotals_112; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_114;
  reg [12:0] frequencyTotals_113; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_115;
  reg [12:0] frequencyTotals_114; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_116;
  reg [12:0] frequencyTotals_115; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_117;
  reg [12:0] frequencyTotals_116; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_118;
  reg [12:0] frequencyTotals_117; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_119;
  reg [12:0] frequencyTotals_118; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_120;
  reg [12:0] frequencyTotals_119; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_121;
  reg [12:0] frequencyTotals_120; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_122;
  reg [12:0] frequencyTotals_121; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_123;
  reg [12:0] frequencyTotals_122; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_124;
  reg [12:0] frequencyTotals_123; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_125;
  reg [12:0] frequencyTotals_124; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_126;
  reg [12:0] frequencyTotals_125; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_127;
  reg [12:0] frequencyTotals_126; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_128;
  reg [12:0] frequencyTotals_127; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_129;
  reg [12:0] frequencyTotals_128; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_130;
  reg [12:0] frequencyTotals_129; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_131;
  reg [12:0] frequencyTotals_130; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_132;
  reg [12:0] frequencyTotals_131; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_133;
  reg [12:0] frequencyTotals_132; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_134;
  reg [12:0] frequencyTotals_133; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_135;
  reg [12:0] frequencyTotals_134; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_136;
  reg [12:0] frequencyTotals_135; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_137;
  reg [12:0] frequencyTotals_136; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_138;
  reg [12:0] frequencyTotals_137; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_139;
  reg [12:0] frequencyTotals_138; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_140;
  reg [12:0] frequencyTotals_139; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_141;
  reg [12:0] frequencyTotals_140; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_142;
  reg [12:0] frequencyTotals_141; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_143;
  reg [12:0] frequencyTotals_142; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_144;
  reg [12:0] frequencyTotals_143; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_145;
  reg [12:0] frequencyTotals_144; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_146;
  reg [12:0] frequencyTotals_145; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_147;
  reg [12:0] frequencyTotals_146; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_148;
  reg [12:0] frequencyTotals_147; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_149;
  reg [12:0] frequencyTotals_148; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_150;
  reg [12:0] frequencyTotals_149; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_151;
  reg [12:0] frequencyTotals_150; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_152;
  reg [12:0] frequencyTotals_151; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_153;
  reg [12:0] frequencyTotals_152; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_154;
  reg [12:0] frequencyTotals_153; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_155;
  reg [12:0] frequencyTotals_154; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_156;
  reg [12:0] frequencyTotals_155; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_157;
  reg [12:0] frequencyTotals_156; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_158;
  reg [12:0] frequencyTotals_157; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_159;
  reg [12:0] frequencyTotals_158; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_160;
  reg [12:0] frequencyTotals_159; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_161;
  reg [12:0] frequencyTotals_160; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_162;
  reg [12:0] frequencyTotals_161; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_163;
  reg [12:0] frequencyTotals_162; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_164;
  reg [12:0] frequencyTotals_163; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_165;
  reg [12:0] frequencyTotals_164; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_166;
  reg [12:0] frequencyTotals_165; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_167;
  reg [12:0] frequencyTotals_166; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_168;
  reg [12:0] frequencyTotals_167; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_169;
  reg [12:0] frequencyTotals_168; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_170;
  reg [12:0] frequencyTotals_169; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_171;
  reg [12:0] frequencyTotals_170; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_172;
  reg [12:0] frequencyTotals_171; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_173;
  reg [12:0] frequencyTotals_172; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_174;
  reg [12:0] frequencyTotals_173; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_175;
  reg [12:0] frequencyTotals_174; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_176;
  reg [12:0] frequencyTotals_175; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_177;
  reg [12:0] frequencyTotals_176; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_178;
  reg [12:0] frequencyTotals_177; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_179;
  reg [12:0] frequencyTotals_178; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_180;
  reg [12:0] frequencyTotals_179; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_181;
  reg [12:0] frequencyTotals_180; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_182;
  reg [12:0] frequencyTotals_181; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_183;
  reg [12:0] frequencyTotals_182; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_184;
  reg [12:0] frequencyTotals_183; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_185;
  reg [12:0] frequencyTotals_184; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_186;
  reg [12:0] frequencyTotals_185; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_187;
  reg [12:0] frequencyTotals_186; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_188;
  reg [12:0] frequencyTotals_187; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_189;
  reg [12:0] frequencyTotals_188; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_190;
  reg [12:0] frequencyTotals_189; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_191;
  reg [12:0] frequencyTotals_190; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_192;
  reg [12:0] frequencyTotals_191; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_193;
  reg [12:0] frequencyTotals_192; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_194;
  reg [12:0] frequencyTotals_193; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_195;
  reg [12:0] frequencyTotals_194; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_196;
  reg [12:0] frequencyTotals_195; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_197;
  reg [12:0] frequencyTotals_196; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_198;
  reg [12:0] frequencyTotals_197; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_199;
  reg [12:0] frequencyTotals_198; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_200;
  reg [12:0] frequencyTotals_199; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_201;
  reg [12:0] frequencyTotals_200; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_202;
  reg [12:0] frequencyTotals_201; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_203;
  reg [12:0] frequencyTotals_202; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_204;
  reg [12:0] frequencyTotals_203; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_205;
  reg [12:0] frequencyTotals_204; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_206;
  reg [12:0] frequencyTotals_205; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_207;
  reg [12:0] frequencyTotals_206; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_208;
  reg [12:0] frequencyTotals_207; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_209;
  reg [12:0] frequencyTotals_208; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_210;
  reg [12:0] frequencyTotals_209; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_211;
  reg [12:0] frequencyTotals_210; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_212;
  reg [12:0] frequencyTotals_211; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_213;
  reg [12:0] frequencyTotals_212; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_214;
  reg [12:0] frequencyTotals_213; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_215;
  reg [12:0] frequencyTotals_214; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_216;
  reg [12:0] frequencyTotals_215; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_217;
  reg [12:0] frequencyTotals_216; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_218;
  reg [12:0] frequencyTotals_217; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_219;
  reg [12:0] frequencyTotals_218; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_220;
  reg [12:0] frequencyTotals_219; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_221;
  reg [12:0] frequencyTotals_220; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_222;
  reg [12:0] frequencyTotals_221; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_223;
  reg [12:0] frequencyTotals_222; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_224;
  reg [12:0] frequencyTotals_223; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_225;
  reg [12:0] frequencyTotals_224; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_226;
  reg [12:0] frequencyTotals_225; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_227;
  reg [12:0] frequencyTotals_226; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_228;
  reg [12:0] frequencyTotals_227; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_229;
  reg [12:0] frequencyTotals_228; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_230;
  reg [12:0] frequencyTotals_229; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_231;
  reg [12:0] frequencyTotals_230; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_232;
  reg [12:0] frequencyTotals_231; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_233;
  reg [12:0] frequencyTotals_232; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_234;
  reg [12:0] frequencyTotals_233; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_235;
  reg [12:0] frequencyTotals_234; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_236;
  reg [12:0] frequencyTotals_235; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_237;
  reg [12:0] frequencyTotals_236; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_238;
  reg [12:0] frequencyTotals_237; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_239;
  reg [12:0] frequencyTotals_238; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_240;
  reg [12:0] frequencyTotals_239; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_241;
  reg [12:0] frequencyTotals_240; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_242;
  reg [12:0] frequencyTotals_241; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_243;
  reg [12:0] frequencyTotals_242; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_244;
  reg [12:0] frequencyTotals_243; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_245;
  reg [12:0] frequencyTotals_244; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_246;
  reg [12:0] frequencyTotals_245; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_247;
  reg [12:0] frequencyTotals_246; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_248;
  reg [12:0] frequencyTotals_247; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_249;
  reg [12:0] frequencyTotals_248; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_250;
  reg [12:0] frequencyTotals_249; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_251;
  reg [12:0] frequencyTotals_250; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_252;
  reg [12:0] frequencyTotals_251; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_253;
  reg [12:0] frequencyTotals_252; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_254;
  reg [12:0] frequencyTotals_253; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_255;
  reg [12:0] frequencyTotals_254; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_256;
  reg [12:0] frequencyTotals_255; // @[characterFrequencyCounter.scala 35:28]
  reg [31:0] _RAND_257;
  wire  _T = ~state; // @[Conditional.scala 37:30]
  wire  _GEN_1 = io_start | state; // @[characterFrequencyCounter.scala 41:22]
  wire  _T_3 = io_dataIn_bits_0 == 8'h0; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1033 = {{12'd0}, _T_3}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_5 = frequencyTotals_0 + _GEN_1033; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_6 = io_dataIn_bits_0 == 8'h1; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1034 = {{12'd0}, _T_6}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_8 = frequencyTotals_1 + _GEN_1034; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_9 = io_dataIn_bits_0 == 8'h2; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1035 = {{12'd0}, _T_9}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_11 = frequencyTotals_2 + _GEN_1035; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_12 = io_dataIn_bits_0 == 8'h3; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1036 = {{12'd0}, _T_12}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_14 = frequencyTotals_3 + _GEN_1036; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_15 = io_dataIn_bits_0 == 8'h4; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1037 = {{12'd0}, _T_15}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_17 = frequencyTotals_4 + _GEN_1037; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_18 = io_dataIn_bits_0 == 8'h5; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1038 = {{12'd0}, _T_18}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_20 = frequencyTotals_5 + _GEN_1038; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_21 = io_dataIn_bits_0 == 8'h6; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1039 = {{12'd0}, _T_21}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_23 = frequencyTotals_6 + _GEN_1039; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_24 = io_dataIn_bits_0 == 8'h7; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1040 = {{12'd0}, _T_24}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_26 = frequencyTotals_7 + _GEN_1040; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_27 = io_dataIn_bits_0 == 8'h8; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1041 = {{12'd0}, _T_27}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_29 = frequencyTotals_8 + _GEN_1041; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_30 = io_dataIn_bits_0 == 8'h9; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1042 = {{12'd0}, _T_30}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_32 = frequencyTotals_9 + _GEN_1042; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_33 = io_dataIn_bits_0 == 8'ha; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1043 = {{12'd0}, _T_33}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_35 = frequencyTotals_10 + _GEN_1043; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_36 = io_dataIn_bits_0 == 8'hb; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1044 = {{12'd0}, _T_36}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_38 = frequencyTotals_11 + _GEN_1044; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_39 = io_dataIn_bits_0 == 8'hc; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1045 = {{12'd0}, _T_39}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_41 = frequencyTotals_12 + _GEN_1045; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_42 = io_dataIn_bits_0 == 8'hd; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1046 = {{12'd0}, _T_42}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_44 = frequencyTotals_13 + _GEN_1046; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_45 = io_dataIn_bits_0 == 8'he; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1047 = {{12'd0}, _T_45}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_47 = frequencyTotals_14 + _GEN_1047; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_48 = io_dataIn_bits_0 == 8'hf; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1048 = {{12'd0}, _T_48}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_50 = frequencyTotals_15 + _GEN_1048; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_51 = io_dataIn_bits_0 == 8'h10; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1049 = {{12'd0}, _T_51}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_53 = frequencyTotals_16 + _GEN_1049; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_54 = io_dataIn_bits_0 == 8'h11; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1050 = {{12'd0}, _T_54}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_56 = frequencyTotals_17 + _GEN_1050; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_57 = io_dataIn_bits_0 == 8'h12; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1051 = {{12'd0}, _T_57}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_59 = frequencyTotals_18 + _GEN_1051; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_60 = io_dataIn_bits_0 == 8'h13; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1052 = {{12'd0}, _T_60}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_62 = frequencyTotals_19 + _GEN_1052; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_63 = io_dataIn_bits_0 == 8'h14; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1053 = {{12'd0}, _T_63}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_65 = frequencyTotals_20 + _GEN_1053; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_66 = io_dataIn_bits_0 == 8'h15; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1054 = {{12'd0}, _T_66}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_68 = frequencyTotals_21 + _GEN_1054; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_69 = io_dataIn_bits_0 == 8'h16; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1055 = {{12'd0}, _T_69}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_71 = frequencyTotals_22 + _GEN_1055; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_72 = io_dataIn_bits_0 == 8'h17; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1056 = {{12'd0}, _T_72}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_74 = frequencyTotals_23 + _GEN_1056; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_75 = io_dataIn_bits_0 == 8'h18; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1057 = {{12'd0}, _T_75}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_77 = frequencyTotals_24 + _GEN_1057; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_78 = io_dataIn_bits_0 == 8'h19; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1058 = {{12'd0}, _T_78}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_80 = frequencyTotals_25 + _GEN_1058; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_81 = io_dataIn_bits_0 == 8'h1a; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1059 = {{12'd0}, _T_81}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_83 = frequencyTotals_26 + _GEN_1059; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_84 = io_dataIn_bits_0 == 8'h1b; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1060 = {{12'd0}, _T_84}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_86 = frequencyTotals_27 + _GEN_1060; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_87 = io_dataIn_bits_0 == 8'h1c; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1061 = {{12'd0}, _T_87}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_89 = frequencyTotals_28 + _GEN_1061; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_90 = io_dataIn_bits_0 == 8'h1d; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1062 = {{12'd0}, _T_90}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_92 = frequencyTotals_29 + _GEN_1062; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_93 = io_dataIn_bits_0 == 8'h1e; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1063 = {{12'd0}, _T_93}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_95 = frequencyTotals_30 + _GEN_1063; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_96 = io_dataIn_bits_0 == 8'h1f; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1064 = {{12'd0}, _T_96}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_98 = frequencyTotals_31 + _GEN_1064; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_99 = io_dataIn_bits_0 == 8'h20; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1065 = {{12'd0}, _T_99}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_101 = frequencyTotals_32 + _GEN_1065; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_102 = io_dataIn_bits_0 == 8'h21; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1066 = {{12'd0}, _T_102}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_104 = frequencyTotals_33 + _GEN_1066; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_105 = io_dataIn_bits_0 == 8'h22; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1067 = {{12'd0}, _T_105}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_107 = frequencyTotals_34 + _GEN_1067; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_108 = io_dataIn_bits_0 == 8'h23; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1068 = {{12'd0}, _T_108}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_110 = frequencyTotals_35 + _GEN_1068; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_111 = io_dataIn_bits_0 == 8'h24; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1069 = {{12'd0}, _T_111}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_113 = frequencyTotals_36 + _GEN_1069; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_114 = io_dataIn_bits_0 == 8'h25; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1070 = {{12'd0}, _T_114}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_116 = frequencyTotals_37 + _GEN_1070; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_117 = io_dataIn_bits_0 == 8'h26; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1071 = {{12'd0}, _T_117}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_119 = frequencyTotals_38 + _GEN_1071; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_120 = io_dataIn_bits_0 == 8'h27; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1072 = {{12'd0}, _T_120}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_122 = frequencyTotals_39 + _GEN_1072; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_123 = io_dataIn_bits_0 == 8'h28; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1073 = {{12'd0}, _T_123}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_125 = frequencyTotals_40 + _GEN_1073; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_126 = io_dataIn_bits_0 == 8'h29; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1074 = {{12'd0}, _T_126}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_128 = frequencyTotals_41 + _GEN_1074; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_129 = io_dataIn_bits_0 == 8'h2a; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1075 = {{12'd0}, _T_129}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_131 = frequencyTotals_42 + _GEN_1075; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_132 = io_dataIn_bits_0 == 8'h2b; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1076 = {{12'd0}, _T_132}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_134 = frequencyTotals_43 + _GEN_1076; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_135 = io_dataIn_bits_0 == 8'h2c; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1077 = {{12'd0}, _T_135}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_137 = frequencyTotals_44 + _GEN_1077; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_138 = io_dataIn_bits_0 == 8'h2d; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1078 = {{12'd0}, _T_138}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_140 = frequencyTotals_45 + _GEN_1078; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_141 = io_dataIn_bits_0 == 8'h2e; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1079 = {{12'd0}, _T_141}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_143 = frequencyTotals_46 + _GEN_1079; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_144 = io_dataIn_bits_0 == 8'h2f; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1080 = {{12'd0}, _T_144}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_146 = frequencyTotals_47 + _GEN_1080; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_147 = io_dataIn_bits_0 == 8'h30; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1081 = {{12'd0}, _T_147}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_149 = frequencyTotals_48 + _GEN_1081; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_150 = io_dataIn_bits_0 == 8'h31; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1082 = {{12'd0}, _T_150}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_152 = frequencyTotals_49 + _GEN_1082; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_153 = io_dataIn_bits_0 == 8'h32; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1083 = {{12'd0}, _T_153}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_155 = frequencyTotals_50 + _GEN_1083; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_156 = io_dataIn_bits_0 == 8'h33; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1084 = {{12'd0}, _T_156}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_158 = frequencyTotals_51 + _GEN_1084; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_159 = io_dataIn_bits_0 == 8'h34; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1085 = {{12'd0}, _T_159}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_161 = frequencyTotals_52 + _GEN_1085; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_162 = io_dataIn_bits_0 == 8'h35; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1086 = {{12'd0}, _T_162}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_164 = frequencyTotals_53 + _GEN_1086; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_165 = io_dataIn_bits_0 == 8'h36; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1087 = {{12'd0}, _T_165}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_167 = frequencyTotals_54 + _GEN_1087; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_168 = io_dataIn_bits_0 == 8'h37; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1088 = {{12'd0}, _T_168}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_170 = frequencyTotals_55 + _GEN_1088; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_171 = io_dataIn_bits_0 == 8'h38; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1089 = {{12'd0}, _T_171}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_173 = frequencyTotals_56 + _GEN_1089; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_174 = io_dataIn_bits_0 == 8'h39; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1090 = {{12'd0}, _T_174}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_176 = frequencyTotals_57 + _GEN_1090; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_177 = io_dataIn_bits_0 == 8'h3a; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1091 = {{12'd0}, _T_177}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_179 = frequencyTotals_58 + _GEN_1091; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_180 = io_dataIn_bits_0 == 8'h3b; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1092 = {{12'd0}, _T_180}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_182 = frequencyTotals_59 + _GEN_1092; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_183 = io_dataIn_bits_0 == 8'h3c; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1093 = {{12'd0}, _T_183}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_185 = frequencyTotals_60 + _GEN_1093; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_186 = io_dataIn_bits_0 == 8'h3d; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1094 = {{12'd0}, _T_186}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_188 = frequencyTotals_61 + _GEN_1094; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_189 = io_dataIn_bits_0 == 8'h3e; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1095 = {{12'd0}, _T_189}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_191 = frequencyTotals_62 + _GEN_1095; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_192 = io_dataIn_bits_0 == 8'h3f; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1096 = {{12'd0}, _T_192}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_194 = frequencyTotals_63 + _GEN_1096; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_195 = io_dataIn_bits_0 == 8'h40; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1097 = {{12'd0}, _T_195}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_197 = frequencyTotals_64 + _GEN_1097; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_198 = io_dataIn_bits_0 == 8'h41; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1098 = {{12'd0}, _T_198}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_200 = frequencyTotals_65 + _GEN_1098; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_201 = io_dataIn_bits_0 == 8'h42; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1099 = {{12'd0}, _T_201}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_203 = frequencyTotals_66 + _GEN_1099; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_204 = io_dataIn_bits_0 == 8'h43; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1100 = {{12'd0}, _T_204}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_206 = frequencyTotals_67 + _GEN_1100; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_207 = io_dataIn_bits_0 == 8'h44; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1101 = {{12'd0}, _T_207}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_209 = frequencyTotals_68 + _GEN_1101; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_210 = io_dataIn_bits_0 == 8'h45; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1102 = {{12'd0}, _T_210}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_212 = frequencyTotals_69 + _GEN_1102; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_213 = io_dataIn_bits_0 == 8'h46; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1103 = {{12'd0}, _T_213}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_215 = frequencyTotals_70 + _GEN_1103; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_216 = io_dataIn_bits_0 == 8'h47; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1104 = {{12'd0}, _T_216}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_218 = frequencyTotals_71 + _GEN_1104; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_219 = io_dataIn_bits_0 == 8'h48; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1105 = {{12'd0}, _T_219}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_221 = frequencyTotals_72 + _GEN_1105; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_222 = io_dataIn_bits_0 == 8'h49; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1106 = {{12'd0}, _T_222}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_224 = frequencyTotals_73 + _GEN_1106; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_225 = io_dataIn_bits_0 == 8'h4a; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1107 = {{12'd0}, _T_225}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_227 = frequencyTotals_74 + _GEN_1107; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_228 = io_dataIn_bits_0 == 8'h4b; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1108 = {{12'd0}, _T_228}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_230 = frequencyTotals_75 + _GEN_1108; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_231 = io_dataIn_bits_0 == 8'h4c; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1109 = {{12'd0}, _T_231}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_233 = frequencyTotals_76 + _GEN_1109; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_234 = io_dataIn_bits_0 == 8'h4d; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1110 = {{12'd0}, _T_234}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_236 = frequencyTotals_77 + _GEN_1110; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_237 = io_dataIn_bits_0 == 8'h4e; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1111 = {{12'd0}, _T_237}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_239 = frequencyTotals_78 + _GEN_1111; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_240 = io_dataIn_bits_0 == 8'h4f; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1112 = {{12'd0}, _T_240}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_242 = frequencyTotals_79 + _GEN_1112; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_243 = io_dataIn_bits_0 == 8'h50; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1113 = {{12'd0}, _T_243}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_245 = frequencyTotals_80 + _GEN_1113; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_246 = io_dataIn_bits_0 == 8'h51; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1114 = {{12'd0}, _T_246}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_248 = frequencyTotals_81 + _GEN_1114; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_249 = io_dataIn_bits_0 == 8'h52; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1115 = {{12'd0}, _T_249}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_251 = frequencyTotals_82 + _GEN_1115; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_252 = io_dataIn_bits_0 == 8'h53; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1116 = {{12'd0}, _T_252}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_254 = frequencyTotals_83 + _GEN_1116; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_255 = io_dataIn_bits_0 == 8'h54; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1117 = {{12'd0}, _T_255}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_257 = frequencyTotals_84 + _GEN_1117; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_258 = io_dataIn_bits_0 == 8'h55; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1118 = {{12'd0}, _T_258}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_260 = frequencyTotals_85 + _GEN_1118; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_261 = io_dataIn_bits_0 == 8'h56; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1119 = {{12'd0}, _T_261}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_263 = frequencyTotals_86 + _GEN_1119; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_264 = io_dataIn_bits_0 == 8'h57; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1120 = {{12'd0}, _T_264}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_266 = frequencyTotals_87 + _GEN_1120; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_267 = io_dataIn_bits_0 == 8'h58; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1121 = {{12'd0}, _T_267}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_269 = frequencyTotals_88 + _GEN_1121; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_270 = io_dataIn_bits_0 == 8'h59; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1122 = {{12'd0}, _T_270}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_272 = frequencyTotals_89 + _GEN_1122; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_273 = io_dataIn_bits_0 == 8'h5a; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1123 = {{12'd0}, _T_273}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_275 = frequencyTotals_90 + _GEN_1123; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_276 = io_dataIn_bits_0 == 8'h5b; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1124 = {{12'd0}, _T_276}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_278 = frequencyTotals_91 + _GEN_1124; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_279 = io_dataIn_bits_0 == 8'h5c; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1125 = {{12'd0}, _T_279}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_281 = frequencyTotals_92 + _GEN_1125; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_282 = io_dataIn_bits_0 == 8'h5d; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1126 = {{12'd0}, _T_282}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_284 = frequencyTotals_93 + _GEN_1126; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_285 = io_dataIn_bits_0 == 8'h5e; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1127 = {{12'd0}, _T_285}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_287 = frequencyTotals_94 + _GEN_1127; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_288 = io_dataIn_bits_0 == 8'h5f; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1128 = {{12'd0}, _T_288}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_290 = frequencyTotals_95 + _GEN_1128; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_291 = io_dataIn_bits_0 == 8'h60; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1129 = {{12'd0}, _T_291}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_293 = frequencyTotals_96 + _GEN_1129; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_294 = io_dataIn_bits_0 == 8'h61; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1130 = {{12'd0}, _T_294}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_296 = frequencyTotals_97 + _GEN_1130; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_297 = io_dataIn_bits_0 == 8'h62; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1131 = {{12'd0}, _T_297}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_299 = frequencyTotals_98 + _GEN_1131; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_300 = io_dataIn_bits_0 == 8'h63; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1132 = {{12'd0}, _T_300}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_302 = frequencyTotals_99 + _GEN_1132; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_303 = io_dataIn_bits_0 == 8'h64; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1133 = {{12'd0}, _T_303}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_305 = frequencyTotals_100 + _GEN_1133; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_306 = io_dataIn_bits_0 == 8'h65; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1134 = {{12'd0}, _T_306}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_308 = frequencyTotals_101 + _GEN_1134; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_309 = io_dataIn_bits_0 == 8'h66; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1135 = {{12'd0}, _T_309}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_311 = frequencyTotals_102 + _GEN_1135; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_312 = io_dataIn_bits_0 == 8'h67; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1136 = {{12'd0}, _T_312}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_314 = frequencyTotals_103 + _GEN_1136; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_315 = io_dataIn_bits_0 == 8'h68; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1137 = {{12'd0}, _T_315}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_317 = frequencyTotals_104 + _GEN_1137; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_318 = io_dataIn_bits_0 == 8'h69; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1138 = {{12'd0}, _T_318}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_320 = frequencyTotals_105 + _GEN_1138; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_321 = io_dataIn_bits_0 == 8'h6a; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1139 = {{12'd0}, _T_321}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_323 = frequencyTotals_106 + _GEN_1139; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_324 = io_dataIn_bits_0 == 8'h6b; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1140 = {{12'd0}, _T_324}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_326 = frequencyTotals_107 + _GEN_1140; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_327 = io_dataIn_bits_0 == 8'h6c; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1141 = {{12'd0}, _T_327}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_329 = frequencyTotals_108 + _GEN_1141; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_330 = io_dataIn_bits_0 == 8'h6d; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1142 = {{12'd0}, _T_330}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_332 = frequencyTotals_109 + _GEN_1142; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_333 = io_dataIn_bits_0 == 8'h6e; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1143 = {{12'd0}, _T_333}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_335 = frequencyTotals_110 + _GEN_1143; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_336 = io_dataIn_bits_0 == 8'h6f; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1144 = {{12'd0}, _T_336}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_338 = frequencyTotals_111 + _GEN_1144; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_339 = io_dataIn_bits_0 == 8'h70; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1145 = {{12'd0}, _T_339}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_341 = frequencyTotals_112 + _GEN_1145; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_342 = io_dataIn_bits_0 == 8'h71; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1146 = {{12'd0}, _T_342}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_344 = frequencyTotals_113 + _GEN_1146; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_345 = io_dataIn_bits_0 == 8'h72; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1147 = {{12'd0}, _T_345}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_347 = frequencyTotals_114 + _GEN_1147; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_348 = io_dataIn_bits_0 == 8'h73; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1148 = {{12'd0}, _T_348}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_350 = frequencyTotals_115 + _GEN_1148; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_351 = io_dataIn_bits_0 == 8'h74; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1149 = {{12'd0}, _T_351}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_353 = frequencyTotals_116 + _GEN_1149; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_354 = io_dataIn_bits_0 == 8'h75; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1150 = {{12'd0}, _T_354}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_356 = frequencyTotals_117 + _GEN_1150; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_357 = io_dataIn_bits_0 == 8'h76; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1151 = {{12'd0}, _T_357}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_359 = frequencyTotals_118 + _GEN_1151; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_360 = io_dataIn_bits_0 == 8'h77; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1152 = {{12'd0}, _T_360}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_362 = frequencyTotals_119 + _GEN_1152; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_363 = io_dataIn_bits_0 == 8'h78; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1153 = {{12'd0}, _T_363}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_365 = frequencyTotals_120 + _GEN_1153; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_366 = io_dataIn_bits_0 == 8'h79; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1154 = {{12'd0}, _T_366}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_368 = frequencyTotals_121 + _GEN_1154; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_369 = io_dataIn_bits_0 == 8'h7a; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1155 = {{12'd0}, _T_369}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_371 = frequencyTotals_122 + _GEN_1155; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_372 = io_dataIn_bits_0 == 8'h7b; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1156 = {{12'd0}, _T_372}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_374 = frequencyTotals_123 + _GEN_1156; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_375 = io_dataIn_bits_0 == 8'h7c; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1157 = {{12'd0}, _T_375}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_377 = frequencyTotals_124 + _GEN_1157; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_378 = io_dataIn_bits_0 == 8'h7d; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1158 = {{12'd0}, _T_378}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_380 = frequencyTotals_125 + _GEN_1158; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_381 = io_dataIn_bits_0 == 8'h7e; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1159 = {{12'd0}, _T_381}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_383 = frequencyTotals_126 + _GEN_1159; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_384 = io_dataIn_bits_0 == 8'h7f; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1160 = {{12'd0}, _T_384}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_386 = frequencyTotals_127 + _GEN_1160; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_387 = io_dataIn_bits_0 == 8'h80; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1161 = {{12'd0}, _T_387}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_389 = frequencyTotals_128 + _GEN_1161; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_390 = io_dataIn_bits_0 == 8'h81; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1162 = {{12'd0}, _T_390}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_392 = frequencyTotals_129 + _GEN_1162; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_393 = io_dataIn_bits_0 == 8'h82; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1163 = {{12'd0}, _T_393}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_395 = frequencyTotals_130 + _GEN_1163; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_396 = io_dataIn_bits_0 == 8'h83; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1164 = {{12'd0}, _T_396}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_398 = frequencyTotals_131 + _GEN_1164; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_399 = io_dataIn_bits_0 == 8'h84; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1165 = {{12'd0}, _T_399}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_401 = frequencyTotals_132 + _GEN_1165; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_402 = io_dataIn_bits_0 == 8'h85; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1166 = {{12'd0}, _T_402}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_404 = frequencyTotals_133 + _GEN_1166; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_405 = io_dataIn_bits_0 == 8'h86; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1167 = {{12'd0}, _T_405}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_407 = frequencyTotals_134 + _GEN_1167; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_408 = io_dataIn_bits_0 == 8'h87; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1168 = {{12'd0}, _T_408}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_410 = frequencyTotals_135 + _GEN_1168; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_411 = io_dataIn_bits_0 == 8'h88; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1169 = {{12'd0}, _T_411}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_413 = frequencyTotals_136 + _GEN_1169; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_414 = io_dataIn_bits_0 == 8'h89; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1170 = {{12'd0}, _T_414}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_416 = frequencyTotals_137 + _GEN_1170; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_417 = io_dataIn_bits_0 == 8'h8a; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1171 = {{12'd0}, _T_417}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_419 = frequencyTotals_138 + _GEN_1171; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_420 = io_dataIn_bits_0 == 8'h8b; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1172 = {{12'd0}, _T_420}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_422 = frequencyTotals_139 + _GEN_1172; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_423 = io_dataIn_bits_0 == 8'h8c; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1173 = {{12'd0}, _T_423}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_425 = frequencyTotals_140 + _GEN_1173; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_426 = io_dataIn_bits_0 == 8'h8d; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1174 = {{12'd0}, _T_426}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_428 = frequencyTotals_141 + _GEN_1174; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_429 = io_dataIn_bits_0 == 8'h8e; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1175 = {{12'd0}, _T_429}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_431 = frequencyTotals_142 + _GEN_1175; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_432 = io_dataIn_bits_0 == 8'h8f; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1176 = {{12'd0}, _T_432}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_434 = frequencyTotals_143 + _GEN_1176; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_435 = io_dataIn_bits_0 == 8'h90; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1177 = {{12'd0}, _T_435}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_437 = frequencyTotals_144 + _GEN_1177; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_438 = io_dataIn_bits_0 == 8'h91; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1178 = {{12'd0}, _T_438}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_440 = frequencyTotals_145 + _GEN_1178; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_441 = io_dataIn_bits_0 == 8'h92; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1179 = {{12'd0}, _T_441}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_443 = frequencyTotals_146 + _GEN_1179; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_444 = io_dataIn_bits_0 == 8'h93; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1180 = {{12'd0}, _T_444}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_446 = frequencyTotals_147 + _GEN_1180; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_447 = io_dataIn_bits_0 == 8'h94; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1181 = {{12'd0}, _T_447}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_449 = frequencyTotals_148 + _GEN_1181; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_450 = io_dataIn_bits_0 == 8'h95; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1182 = {{12'd0}, _T_450}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_452 = frequencyTotals_149 + _GEN_1182; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_453 = io_dataIn_bits_0 == 8'h96; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1183 = {{12'd0}, _T_453}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_455 = frequencyTotals_150 + _GEN_1183; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_456 = io_dataIn_bits_0 == 8'h97; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1184 = {{12'd0}, _T_456}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_458 = frequencyTotals_151 + _GEN_1184; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_459 = io_dataIn_bits_0 == 8'h98; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1185 = {{12'd0}, _T_459}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_461 = frequencyTotals_152 + _GEN_1185; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_462 = io_dataIn_bits_0 == 8'h99; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1186 = {{12'd0}, _T_462}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_464 = frequencyTotals_153 + _GEN_1186; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_465 = io_dataIn_bits_0 == 8'h9a; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1187 = {{12'd0}, _T_465}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_467 = frequencyTotals_154 + _GEN_1187; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_468 = io_dataIn_bits_0 == 8'h9b; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1188 = {{12'd0}, _T_468}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_470 = frequencyTotals_155 + _GEN_1188; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_471 = io_dataIn_bits_0 == 8'h9c; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1189 = {{12'd0}, _T_471}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_473 = frequencyTotals_156 + _GEN_1189; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_474 = io_dataIn_bits_0 == 8'h9d; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1190 = {{12'd0}, _T_474}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_476 = frequencyTotals_157 + _GEN_1190; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_477 = io_dataIn_bits_0 == 8'h9e; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1191 = {{12'd0}, _T_477}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_479 = frequencyTotals_158 + _GEN_1191; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_480 = io_dataIn_bits_0 == 8'h9f; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1192 = {{12'd0}, _T_480}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_482 = frequencyTotals_159 + _GEN_1192; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_483 = io_dataIn_bits_0 == 8'ha0; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1193 = {{12'd0}, _T_483}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_485 = frequencyTotals_160 + _GEN_1193; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_486 = io_dataIn_bits_0 == 8'ha1; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1194 = {{12'd0}, _T_486}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_488 = frequencyTotals_161 + _GEN_1194; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_489 = io_dataIn_bits_0 == 8'ha2; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1195 = {{12'd0}, _T_489}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_491 = frequencyTotals_162 + _GEN_1195; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_492 = io_dataIn_bits_0 == 8'ha3; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1196 = {{12'd0}, _T_492}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_494 = frequencyTotals_163 + _GEN_1196; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_495 = io_dataIn_bits_0 == 8'ha4; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1197 = {{12'd0}, _T_495}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_497 = frequencyTotals_164 + _GEN_1197; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_498 = io_dataIn_bits_0 == 8'ha5; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1198 = {{12'd0}, _T_498}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_500 = frequencyTotals_165 + _GEN_1198; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_501 = io_dataIn_bits_0 == 8'ha6; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1199 = {{12'd0}, _T_501}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_503 = frequencyTotals_166 + _GEN_1199; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_504 = io_dataIn_bits_0 == 8'ha7; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1200 = {{12'd0}, _T_504}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_506 = frequencyTotals_167 + _GEN_1200; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_507 = io_dataIn_bits_0 == 8'ha8; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1201 = {{12'd0}, _T_507}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_509 = frequencyTotals_168 + _GEN_1201; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_510 = io_dataIn_bits_0 == 8'ha9; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1202 = {{12'd0}, _T_510}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_512 = frequencyTotals_169 + _GEN_1202; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_513 = io_dataIn_bits_0 == 8'haa; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1203 = {{12'd0}, _T_513}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_515 = frequencyTotals_170 + _GEN_1203; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_516 = io_dataIn_bits_0 == 8'hab; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1204 = {{12'd0}, _T_516}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_518 = frequencyTotals_171 + _GEN_1204; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_519 = io_dataIn_bits_0 == 8'hac; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1205 = {{12'd0}, _T_519}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_521 = frequencyTotals_172 + _GEN_1205; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_522 = io_dataIn_bits_0 == 8'had; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1206 = {{12'd0}, _T_522}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_524 = frequencyTotals_173 + _GEN_1206; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_525 = io_dataIn_bits_0 == 8'hae; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1207 = {{12'd0}, _T_525}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_527 = frequencyTotals_174 + _GEN_1207; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_528 = io_dataIn_bits_0 == 8'haf; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1208 = {{12'd0}, _T_528}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_530 = frequencyTotals_175 + _GEN_1208; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_531 = io_dataIn_bits_0 == 8'hb0; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1209 = {{12'd0}, _T_531}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_533 = frequencyTotals_176 + _GEN_1209; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_534 = io_dataIn_bits_0 == 8'hb1; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1210 = {{12'd0}, _T_534}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_536 = frequencyTotals_177 + _GEN_1210; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_537 = io_dataIn_bits_0 == 8'hb2; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1211 = {{12'd0}, _T_537}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_539 = frequencyTotals_178 + _GEN_1211; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_540 = io_dataIn_bits_0 == 8'hb3; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1212 = {{12'd0}, _T_540}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_542 = frequencyTotals_179 + _GEN_1212; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_543 = io_dataIn_bits_0 == 8'hb4; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1213 = {{12'd0}, _T_543}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_545 = frequencyTotals_180 + _GEN_1213; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_546 = io_dataIn_bits_0 == 8'hb5; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1214 = {{12'd0}, _T_546}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_548 = frequencyTotals_181 + _GEN_1214; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_549 = io_dataIn_bits_0 == 8'hb6; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1215 = {{12'd0}, _T_549}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_551 = frequencyTotals_182 + _GEN_1215; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_552 = io_dataIn_bits_0 == 8'hb7; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1216 = {{12'd0}, _T_552}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_554 = frequencyTotals_183 + _GEN_1216; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_555 = io_dataIn_bits_0 == 8'hb8; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1217 = {{12'd0}, _T_555}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_557 = frequencyTotals_184 + _GEN_1217; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_558 = io_dataIn_bits_0 == 8'hb9; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1218 = {{12'd0}, _T_558}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_560 = frequencyTotals_185 + _GEN_1218; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_561 = io_dataIn_bits_0 == 8'hba; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1219 = {{12'd0}, _T_561}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_563 = frequencyTotals_186 + _GEN_1219; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_564 = io_dataIn_bits_0 == 8'hbb; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1220 = {{12'd0}, _T_564}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_566 = frequencyTotals_187 + _GEN_1220; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_567 = io_dataIn_bits_0 == 8'hbc; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1221 = {{12'd0}, _T_567}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_569 = frequencyTotals_188 + _GEN_1221; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_570 = io_dataIn_bits_0 == 8'hbd; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1222 = {{12'd0}, _T_570}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_572 = frequencyTotals_189 + _GEN_1222; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_573 = io_dataIn_bits_0 == 8'hbe; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1223 = {{12'd0}, _T_573}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_575 = frequencyTotals_190 + _GEN_1223; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_576 = io_dataIn_bits_0 == 8'hbf; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1224 = {{12'd0}, _T_576}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_578 = frequencyTotals_191 + _GEN_1224; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_579 = io_dataIn_bits_0 == 8'hc0; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1225 = {{12'd0}, _T_579}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_581 = frequencyTotals_192 + _GEN_1225; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_582 = io_dataIn_bits_0 == 8'hc1; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1226 = {{12'd0}, _T_582}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_584 = frequencyTotals_193 + _GEN_1226; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_585 = io_dataIn_bits_0 == 8'hc2; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1227 = {{12'd0}, _T_585}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_587 = frequencyTotals_194 + _GEN_1227; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_588 = io_dataIn_bits_0 == 8'hc3; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1228 = {{12'd0}, _T_588}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_590 = frequencyTotals_195 + _GEN_1228; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_591 = io_dataIn_bits_0 == 8'hc4; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1229 = {{12'd0}, _T_591}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_593 = frequencyTotals_196 + _GEN_1229; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_594 = io_dataIn_bits_0 == 8'hc5; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1230 = {{12'd0}, _T_594}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_596 = frequencyTotals_197 + _GEN_1230; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_597 = io_dataIn_bits_0 == 8'hc6; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1231 = {{12'd0}, _T_597}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_599 = frequencyTotals_198 + _GEN_1231; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_600 = io_dataIn_bits_0 == 8'hc7; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1232 = {{12'd0}, _T_600}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_602 = frequencyTotals_199 + _GEN_1232; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_603 = io_dataIn_bits_0 == 8'hc8; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1233 = {{12'd0}, _T_603}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_605 = frequencyTotals_200 + _GEN_1233; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_606 = io_dataIn_bits_0 == 8'hc9; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1234 = {{12'd0}, _T_606}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_608 = frequencyTotals_201 + _GEN_1234; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_609 = io_dataIn_bits_0 == 8'hca; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1235 = {{12'd0}, _T_609}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_611 = frequencyTotals_202 + _GEN_1235; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_612 = io_dataIn_bits_0 == 8'hcb; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1236 = {{12'd0}, _T_612}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_614 = frequencyTotals_203 + _GEN_1236; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_615 = io_dataIn_bits_0 == 8'hcc; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1237 = {{12'd0}, _T_615}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_617 = frequencyTotals_204 + _GEN_1237; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_618 = io_dataIn_bits_0 == 8'hcd; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1238 = {{12'd0}, _T_618}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_620 = frequencyTotals_205 + _GEN_1238; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_621 = io_dataIn_bits_0 == 8'hce; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1239 = {{12'd0}, _T_621}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_623 = frequencyTotals_206 + _GEN_1239; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_624 = io_dataIn_bits_0 == 8'hcf; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1240 = {{12'd0}, _T_624}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_626 = frequencyTotals_207 + _GEN_1240; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_627 = io_dataIn_bits_0 == 8'hd0; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1241 = {{12'd0}, _T_627}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_629 = frequencyTotals_208 + _GEN_1241; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_630 = io_dataIn_bits_0 == 8'hd1; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1242 = {{12'd0}, _T_630}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_632 = frequencyTotals_209 + _GEN_1242; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_633 = io_dataIn_bits_0 == 8'hd2; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1243 = {{12'd0}, _T_633}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_635 = frequencyTotals_210 + _GEN_1243; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_636 = io_dataIn_bits_0 == 8'hd3; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1244 = {{12'd0}, _T_636}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_638 = frequencyTotals_211 + _GEN_1244; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_639 = io_dataIn_bits_0 == 8'hd4; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1245 = {{12'd0}, _T_639}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_641 = frequencyTotals_212 + _GEN_1245; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_642 = io_dataIn_bits_0 == 8'hd5; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1246 = {{12'd0}, _T_642}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_644 = frequencyTotals_213 + _GEN_1246; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_645 = io_dataIn_bits_0 == 8'hd6; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1247 = {{12'd0}, _T_645}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_647 = frequencyTotals_214 + _GEN_1247; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_648 = io_dataIn_bits_0 == 8'hd7; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1248 = {{12'd0}, _T_648}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_650 = frequencyTotals_215 + _GEN_1248; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_651 = io_dataIn_bits_0 == 8'hd8; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1249 = {{12'd0}, _T_651}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_653 = frequencyTotals_216 + _GEN_1249; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_654 = io_dataIn_bits_0 == 8'hd9; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1250 = {{12'd0}, _T_654}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_656 = frequencyTotals_217 + _GEN_1250; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_657 = io_dataIn_bits_0 == 8'hda; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1251 = {{12'd0}, _T_657}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_659 = frequencyTotals_218 + _GEN_1251; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_660 = io_dataIn_bits_0 == 8'hdb; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1252 = {{12'd0}, _T_660}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_662 = frequencyTotals_219 + _GEN_1252; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_663 = io_dataIn_bits_0 == 8'hdc; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1253 = {{12'd0}, _T_663}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_665 = frequencyTotals_220 + _GEN_1253; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_666 = io_dataIn_bits_0 == 8'hdd; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1254 = {{12'd0}, _T_666}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_668 = frequencyTotals_221 + _GEN_1254; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_669 = io_dataIn_bits_0 == 8'hde; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1255 = {{12'd0}, _T_669}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_671 = frequencyTotals_222 + _GEN_1255; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_672 = io_dataIn_bits_0 == 8'hdf; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1256 = {{12'd0}, _T_672}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_674 = frequencyTotals_223 + _GEN_1256; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_675 = io_dataIn_bits_0 == 8'he0; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1257 = {{12'd0}, _T_675}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_677 = frequencyTotals_224 + _GEN_1257; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_678 = io_dataIn_bits_0 == 8'he1; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1258 = {{12'd0}, _T_678}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_680 = frequencyTotals_225 + _GEN_1258; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_681 = io_dataIn_bits_0 == 8'he2; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1259 = {{12'd0}, _T_681}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_683 = frequencyTotals_226 + _GEN_1259; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_684 = io_dataIn_bits_0 == 8'he3; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1260 = {{12'd0}, _T_684}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_686 = frequencyTotals_227 + _GEN_1260; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_687 = io_dataIn_bits_0 == 8'he4; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1261 = {{12'd0}, _T_687}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_689 = frequencyTotals_228 + _GEN_1261; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_690 = io_dataIn_bits_0 == 8'he5; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1262 = {{12'd0}, _T_690}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_692 = frequencyTotals_229 + _GEN_1262; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_693 = io_dataIn_bits_0 == 8'he6; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1263 = {{12'd0}, _T_693}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_695 = frequencyTotals_230 + _GEN_1263; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_696 = io_dataIn_bits_0 == 8'he7; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1264 = {{12'd0}, _T_696}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_698 = frequencyTotals_231 + _GEN_1264; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_699 = io_dataIn_bits_0 == 8'he8; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1265 = {{12'd0}, _T_699}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_701 = frequencyTotals_232 + _GEN_1265; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_702 = io_dataIn_bits_0 == 8'he9; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1266 = {{12'd0}, _T_702}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_704 = frequencyTotals_233 + _GEN_1266; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_705 = io_dataIn_bits_0 == 8'hea; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1267 = {{12'd0}, _T_705}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_707 = frequencyTotals_234 + _GEN_1267; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_708 = io_dataIn_bits_0 == 8'heb; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1268 = {{12'd0}, _T_708}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_710 = frequencyTotals_235 + _GEN_1268; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_711 = io_dataIn_bits_0 == 8'hec; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1269 = {{12'd0}, _T_711}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_713 = frequencyTotals_236 + _GEN_1269; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_714 = io_dataIn_bits_0 == 8'hed; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1270 = {{12'd0}, _T_714}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_716 = frequencyTotals_237 + _GEN_1270; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_717 = io_dataIn_bits_0 == 8'hee; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1271 = {{12'd0}, _T_717}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_719 = frequencyTotals_238 + _GEN_1271; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_720 = io_dataIn_bits_0 == 8'hef; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1272 = {{12'd0}, _T_720}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_722 = frequencyTotals_239 + _GEN_1272; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_723 = io_dataIn_bits_0 == 8'hf0; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1273 = {{12'd0}, _T_723}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_725 = frequencyTotals_240 + _GEN_1273; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_726 = io_dataIn_bits_0 == 8'hf1; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1274 = {{12'd0}, _T_726}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_728 = frequencyTotals_241 + _GEN_1274; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_729 = io_dataIn_bits_0 == 8'hf2; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1275 = {{12'd0}, _T_729}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_731 = frequencyTotals_242 + _GEN_1275; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_732 = io_dataIn_bits_0 == 8'hf3; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1276 = {{12'd0}, _T_732}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_734 = frequencyTotals_243 + _GEN_1276; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_735 = io_dataIn_bits_0 == 8'hf4; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1277 = {{12'd0}, _T_735}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_737 = frequencyTotals_244 + _GEN_1277; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_738 = io_dataIn_bits_0 == 8'hf5; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1278 = {{12'd0}, _T_738}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_740 = frequencyTotals_245 + _GEN_1278; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_741 = io_dataIn_bits_0 == 8'hf6; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1279 = {{12'd0}, _T_741}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_743 = frequencyTotals_246 + _GEN_1279; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_744 = io_dataIn_bits_0 == 8'hf7; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1280 = {{12'd0}, _T_744}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_746 = frequencyTotals_247 + _GEN_1280; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_747 = io_dataIn_bits_0 == 8'hf8; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1281 = {{12'd0}, _T_747}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_749 = frequencyTotals_248 + _GEN_1281; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_750 = io_dataIn_bits_0 == 8'hf9; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1282 = {{12'd0}, _T_750}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_752 = frequencyTotals_249 + _GEN_1282; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_753 = io_dataIn_bits_0 == 8'hfa; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1283 = {{12'd0}, _T_753}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_755 = frequencyTotals_250 + _GEN_1283; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_756 = io_dataIn_bits_0 == 8'hfb; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1284 = {{12'd0}, _T_756}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_758 = frequencyTotals_251 + _GEN_1284; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_759 = io_dataIn_bits_0 == 8'hfc; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1285 = {{12'd0}, _T_759}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_761 = frequencyTotals_252 + _GEN_1285; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_762 = io_dataIn_bits_0 == 8'hfd; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1286 = {{12'd0}, _T_762}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_764 = frequencyTotals_253 + _GEN_1286; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_765 = io_dataIn_bits_0 == 8'hfe; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1287 = {{12'd0}, _T_765}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_767 = frequencyTotals_254 + _GEN_1287; // @[characterFrequencyCounter.scala 57:60]
  wire  _T_768 = io_dataIn_bits_0 == 8'hff; // @[characterFrequencyCounter.scala 58:43]
  wire [12:0] _GEN_1288 = {{12'd0}, _T_768}; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_770 = frequencyTotals_255 + _GEN_1288; // @[characterFrequencyCounter.scala 57:60]
  wire [12:0] _T_772 = currentByte + 13'h1; // @[characterFrequencyCounter.scala 60:36]
  wire  _T_773 = currentByte >= 13'hfff; // @[characterFrequencyCounter.scala 61:26]
  assign io_dataIn_ready = state; // @[characterFrequencyCounter.scala 71:19]
  assign io_currentByte = currentByte[11:0]; // @[characterFrequencyCounter.scala 68:18]
  assign io_frequencies_0 = frequencyTotals_0; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_1 = frequencyTotals_1; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_2 = frequencyTotals_2; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_3 = frequencyTotals_3; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_4 = frequencyTotals_4; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_5 = frequencyTotals_5; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_6 = frequencyTotals_6; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_7 = frequencyTotals_7; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_8 = frequencyTotals_8; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_9 = frequencyTotals_9; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_10 = frequencyTotals_10; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_11 = frequencyTotals_11; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_12 = frequencyTotals_12; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_13 = frequencyTotals_13; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_14 = frequencyTotals_14; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_15 = frequencyTotals_15; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_16 = frequencyTotals_16; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_17 = frequencyTotals_17; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_18 = frequencyTotals_18; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_19 = frequencyTotals_19; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_20 = frequencyTotals_20; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_21 = frequencyTotals_21; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_22 = frequencyTotals_22; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_23 = frequencyTotals_23; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_24 = frequencyTotals_24; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_25 = frequencyTotals_25; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_26 = frequencyTotals_26; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_27 = frequencyTotals_27; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_28 = frequencyTotals_28; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_29 = frequencyTotals_29; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_30 = frequencyTotals_30; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_31 = frequencyTotals_31; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_32 = frequencyTotals_32; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_33 = frequencyTotals_33; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_34 = frequencyTotals_34; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_35 = frequencyTotals_35; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_36 = frequencyTotals_36; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_37 = frequencyTotals_37; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_38 = frequencyTotals_38; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_39 = frequencyTotals_39; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_40 = frequencyTotals_40; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_41 = frequencyTotals_41; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_42 = frequencyTotals_42; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_43 = frequencyTotals_43; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_44 = frequencyTotals_44; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_45 = frequencyTotals_45; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_46 = frequencyTotals_46; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_47 = frequencyTotals_47; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_48 = frequencyTotals_48; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_49 = frequencyTotals_49; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_50 = frequencyTotals_50; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_51 = frequencyTotals_51; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_52 = frequencyTotals_52; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_53 = frequencyTotals_53; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_54 = frequencyTotals_54; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_55 = frequencyTotals_55; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_56 = frequencyTotals_56; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_57 = frequencyTotals_57; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_58 = frequencyTotals_58; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_59 = frequencyTotals_59; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_60 = frequencyTotals_60; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_61 = frequencyTotals_61; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_62 = frequencyTotals_62; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_63 = frequencyTotals_63; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_64 = frequencyTotals_64; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_65 = frequencyTotals_65; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_66 = frequencyTotals_66; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_67 = frequencyTotals_67; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_68 = frequencyTotals_68; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_69 = frequencyTotals_69; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_70 = frequencyTotals_70; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_71 = frequencyTotals_71; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_72 = frequencyTotals_72; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_73 = frequencyTotals_73; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_74 = frequencyTotals_74; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_75 = frequencyTotals_75; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_76 = frequencyTotals_76; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_77 = frequencyTotals_77; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_78 = frequencyTotals_78; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_79 = frequencyTotals_79; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_80 = frequencyTotals_80; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_81 = frequencyTotals_81; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_82 = frequencyTotals_82; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_83 = frequencyTotals_83; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_84 = frequencyTotals_84; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_85 = frequencyTotals_85; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_86 = frequencyTotals_86; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_87 = frequencyTotals_87; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_88 = frequencyTotals_88; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_89 = frequencyTotals_89; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_90 = frequencyTotals_90; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_91 = frequencyTotals_91; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_92 = frequencyTotals_92; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_93 = frequencyTotals_93; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_94 = frequencyTotals_94; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_95 = frequencyTotals_95; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_96 = frequencyTotals_96; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_97 = frequencyTotals_97; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_98 = frequencyTotals_98; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_99 = frequencyTotals_99; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_100 = frequencyTotals_100; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_101 = frequencyTotals_101; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_102 = frequencyTotals_102; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_103 = frequencyTotals_103; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_104 = frequencyTotals_104; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_105 = frequencyTotals_105; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_106 = frequencyTotals_106; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_107 = frequencyTotals_107; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_108 = frequencyTotals_108; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_109 = frequencyTotals_109; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_110 = frequencyTotals_110; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_111 = frequencyTotals_111; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_112 = frequencyTotals_112; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_113 = frequencyTotals_113; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_114 = frequencyTotals_114; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_115 = frequencyTotals_115; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_116 = frequencyTotals_116; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_117 = frequencyTotals_117; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_118 = frequencyTotals_118; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_119 = frequencyTotals_119; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_120 = frequencyTotals_120; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_121 = frequencyTotals_121; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_122 = frequencyTotals_122; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_123 = frequencyTotals_123; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_124 = frequencyTotals_124; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_125 = frequencyTotals_125; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_126 = frequencyTotals_126; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_127 = frequencyTotals_127; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_128 = frequencyTotals_128; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_129 = frequencyTotals_129; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_130 = frequencyTotals_130; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_131 = frequencyTotals_131; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_132 = frequencyTotals_132; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_133 = frequencyTotals_133; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_134 = frequencyTotals_134; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_135 = frequencyTotals_135; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_136 = frequencyTotals_136; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_137 = frequencyTotals_137; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_138 = frequencyTotals_138; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_139 = frequencyTotals_139; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_140 = frequencyTotals_140; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_141 = frequencyTotals_141; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_142 = frequencyTotals_142; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_143 = frequencyTotals_143; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_144 = frequencyTotals_144; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_145 = frequencyTotals_145; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_146 = frequencyTotals_146; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_147 = frequencyTotals_147; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_148 = frequencyTotals_148; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_149 = frequencyTotals_149; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_150 = frequencyTotals_150; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_151 = frequencyTotals_151; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_152 = frequencyTotals_152; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_153 = frequencyTotals_153; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_154 = frequencyTotals_154; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_155 = frequencyTotals_155; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_156 = frequencyTotals_156; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_157 = frequencyTotals_157; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_158 = frequencyTotals_158; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_159 = frequencyTotals_159; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_160 = frequencyTotals_160; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_161 = frequencyTotals_161; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_162 = frequencyTotals_162; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_163 = frequencyTotals_163; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_164 = frequencyTotals_164; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_165 = frequencyTotals_165; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_166 = frequencyTotals_166; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_167 = frequencyTotals_167; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_168 = frequencyTotals_168; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_169 = frequencyTotals_169; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_170 = frequencyTotals_170; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_171 = frequencyTotals_171; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_172 = frequencyTotals_172; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_173 = frequencyTotals_173; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_174 = frequencyTotals_174; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_175 = frequencyTotals_175; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_176 = frequencyTotals_176; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_177 = frequencyTotals_177; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_178 = frequencyTotals_178; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_179 = frequencyTotals_179; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_180 = frequencyTotals_180; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_181 = frequencyTotals_181; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_182 = frequencyTotals_182; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_183 = frequencyTotals_183; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_184 = frequencyTotals_184; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_185 = frequencyTotals_185; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_186 = frequencyTotals_186; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_187 = frequencyTotals_187; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_188 = frequencyTotals_188; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_189 = frequencyTotals_189; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_190 = frequencyTotals_190; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_191 = frequencyTotals_191; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_192 = frequencyTotals_192; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_193 = frequencyTotals_193; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_194 = frequencyTotals_194; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_195 = frequencyTotals_195; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_196 = frequencyTotals_196; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_197 = frequencyTotals_197; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_198 = frequencyTotals_198; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_199 = frequencyTotals_199; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_200 = frequencyTotals_200; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_201 = frequencyTotals_201; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_202 = frequencyTotals_202; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_203 = frequencyTotals_203; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_204 = frequencyTotals_204; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_205 = frequencyTotals_205; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_206 = frequencyTotals_206; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_207 = frequencyTotals_207; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_208 = frequencyTotals_208; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_209 = frequencyTotals_209; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_210 = frequencyTotals_210; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_211 = frequencyTotals_211; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_212 = frequencyTotals_212; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_213 = frequencyTotals_213; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_214 = frequencyTotals_214; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_215 = frequencyTotals_215; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_216 = frequencyTotals_216; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_217 = frequencyTotals_217; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_218 = frequencyTotals_218; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_219 = frequencyTotals_219; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_220 = frequencyTotals_220; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_221 = frequencyTotals_221; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_222 = frequencyTotals_222; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_223 = frequencyTotals_223; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_224 = frequencyTotals_224; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_225 = frequencyTotals_225; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_226 = frequencyTotals_226; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_227 = frequencyTotals_227; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_228 = frequencyTotals_228; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_229 = frequencyTotals_229; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_230 = frequencyTotals_230; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_231 = frequencyTotals_231; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_232 = frequencyTotals_232; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_233 = frequencyTotals_233; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_234 = frequencyTotals_234; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_235 = frequencyTotals_235; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_236 = frequencyTotals_236; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_237 = frequencyTotals_237; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_238 = frequencyTotals_238; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_239 = frequencyTotals_239; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_240 = frequencyTotals_240; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_241 = frequencyTotals_241; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_242 = frequencyTotals_242; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_243 = frequencyTotals_243; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_244 = frequencyTotals_244; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_245 = frequencyTotals_245; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_246 = frequencyTotals_246; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_247 = frequencyTotals_247; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_248 = frequencyTotals_248; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_249 = frequencyTotals_249; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_250 = frequencyTotals_250; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_251 = frequencyTotals_251; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_252 = frequencyTotals_252; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_253 = frequencyTotals_253; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_254 = frequencyTotals_254; // @[characterFrequencyCounter.scala 69:18]
  assign io_frequencies_255 = frequencyTotals_255; // @[characterFrequencyCounter.scala 69:18]
  assign io_finished = ~state; // @[characterFrequencyCounter.scala 70:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  currentByte = _RAND_1[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  frequencyTotals_0 = _RAND_2[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  frequencyTotals_1 = _RAND_3[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  frequencyTotals_2 = _RAND_4[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  frequencyTotals_3 = _RAND_5[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  frequencyTotals_4 = _RAND_6[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  frequencyTotals_5 = _RAND_7[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  frequencyTotals_6 = _RAND_8[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  frequencyTotals_7 = _RAND_9[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  frequencyTotals_8 = _RAND_10[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  frequencyTotals_9 = _RAND_11[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  frequencyTotals_10 = _RAND_12[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  frequencyTotals_11 = _RAND_13[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  frequencyTotals_12 = _RAND_14[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  frequencyTotals_13 = _RAND_15[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  frequencyTotals_14 = _RAND_16[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  frequencyTotals_15 = _RAND_17[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  frequencyTotals_16 = _RAND_18[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  frequencyTotals_17 = _RAND_19[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  frequencyTotals_18 = _RAND_20[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  frequencyTotals_19 = _RAND_21[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  frequencyTotals_20 = _RAND_22[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  frequencyTotals_21 = _RAND_23[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  frequencyTotals_22 = _RAND_24[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  frequencyTotals_23 = _RAND_25[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  frequencyTotals_24 = _RAND_26[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  frequencyTotals_25 = _RAND_27[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  frequencyTotals_26 = _RAND_28[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  frequencyTotals_27 = _RAND_29[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  frequencyTotals_28 = _RAND_30[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  frequencyTotals_29 = _RAND_31[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  frequencyTotals_30 = _RAND_32[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  frequencyTotals_31 = _RAND_33[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  frequencyTotals_32 = _RAND_34[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  frequencyTotals_33 = _RAND_35[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  frequencyTotals_34 = _RAND_36[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  frequencyTotals_35 = _RAND_37[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  frequencyTotals_36 = _RAND_38[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  frequencyTotals_37 = _RAND_39[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  frequencyTotals_38 = _RAND_40[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  frequencyTotals_39 = _RAND_41[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  frequencyTotals_40 = _RAND_42[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  frequencyTotals_41 = _RAND_43[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  frequencyTotals_42 = _RAND_44[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  frequencyTotals_43 = _RAND_45[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  frequencyTotals_44 = _RAND_46[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  frequencyTotals_45 = _RAND_47[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  frequencyTotals_46 = _RAND_48[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  frequencyTotals_47 = _RAND_49[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  frequencyTotals_48 = _RAND_50[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  frequencyTotals_49 = _RAND_51[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  frequencyTotals_50 = _RAND_52[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  frequencyTotals_51 = _RAND_53[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  frequencyTotals_52 = _RAND_54[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  frequencyTotals_53 = _RAND_55[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  frequencyTotals_54 = _RAND_56[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  frequencyTotals_55 = _RAND_57[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  frequencyTotals_56 = _RAND_58[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  frequencyTotals_57 = _RAND_59[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  frequencyTotals_58 = _RAND_60[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  frequencyTotals_59 = _RAND_61[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  frequencyTotals_60 = _RAND_62[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  frequencyTotals_61 = _RAND_63[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  frequencyTotals_62 = _RAND_64[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  frequencyTotals_63 = _RAND_65[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  frequencyTotals_64 = _RAND_66[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  frequencyTotals_65 = _RAND_67[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  frequencyTotals_66 = _RAND_68[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  frequencyTotals_67 = _RAND_69[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  frequencyTotals_68 = _RAND_70[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  frequencyTotals_69 = _RAND_71[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  frequencyTotals_70 = _RAND_72[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  frequencyTotals_71 = _RAND_73[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  frequencyTotals_72 = _RAND_74[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  frequencyTotals_73 = _RAND_75[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  frequencyTotals_74 = _RAND_76[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  frequencyTotals_75 = _RAND_77[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  frequencyTotals_76 = _RAND_78[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  frequencyTotals_77 = _RAND_79[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  frequencyTotals_78 = _RAND_80[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  frequencyTotals_79 = _RAND_81[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  frequencyTotals_80 = _RAND_82[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  frequencyTotals_81 = _RAND_83[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  frequencyTotals_82 = _RAND_84[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  frequencyTotals_83 = _RAND_85[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  frequencyTotals_84 = _RAND_86[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  frequencyTotals_85 = _RAND_87[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  frequencyTotals_86 = _RAND_88[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  frequencyTotals_87 = _RAND_89[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  frequencyTotals_88 = _RAND_90[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  frequencyTotals_89 = _RAND_91[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  frequencyTotals_90 = _RAND_92[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  frequencyTotals_91 = _RAND_93[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  frequencyTotals_92 = _RAND_94[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  frequencyTotals_93 = _RAND_95[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  frequencyTotals_94 = _RAND_96[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  frequencyTotals_95 = _RAND_97[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  frequencyTotals_96 = _RAND_98[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  frequencyTotals_97 = _RAND_99[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  frequencyTotals_98 = _RAND_100[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  frequencyTotals_99 = _RAND_101[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  frequencyTotals_100 = _RAND_102[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  frequencyTotals_101 = _RAND_103[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  frequencyTotals_102 = _RAND_104[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  frequencyTotals_103 = _RAND_105[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  frequencyTotals_104 = _RAND_106[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  frequencyTotals_105 = _RAND_107[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  frequencyTotals_106 = _RAND_108[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  frequencyTotals_107 = _RAND_109[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  frequencyTotals_108 = _RAND_110[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  frequencyTotals_109 = _RAND_111[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  frequencyTotals_110 = _RAND_112[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  frequencyTotals_111 = _RAND_113[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  frequencyTotals_112 = _RAND_114[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  frequencyTotals_113 = _RAND_115[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  frequencyTotals_114 = _RAND_116[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  frequencyTotals_115 = _RAND_117[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  frequencyTotals_116 = _RAND_118[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  frequencyTotals_117 = _RAND_119[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  frequencyTotals_118 = _RAND_120[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  frequencyTotals_119 = _RAND_121[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  frequencyTotals_120 = _RAND_122[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  frequencyTotals_121 = _RAND_123[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  frequencyTotals_122 = _RAND_124[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  frequencyTotals_123 = _RAND_125[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  frequencyTotals_124 = _RAND_126[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  frequencyTotals_125 = _RAND_127[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  frequencyTotals_126 = _RAND_128[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  frequencyTotals_127 = _RAND_129[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  frequencyTotals_128 = _RAND_130[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  frequencyTotals_129 = _RAND_131[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  frequencyTotals_130 = _RAND_132[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  frequencyTotals_131 = _RAND_133[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  frequencyTotals_132 = _RAND_134[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  frequencyTotals_133 = _RAND_135[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  frequencyTotals_134 = _RAND_136[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  frequencyTotals_135 = _RAND_137[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  frequencyTotals_136 = _RAND_138[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  frequencyTotals_137 = _RAND_139[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  frequencyTotals_138 = _RAND_140[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  frequencyTotals_139 = _RAND_141[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  frequencyTotals_140 = _RAND_142[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  frequencyTotals_141 = _RAND_143[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  frequencyTotals_142 = _RAND_144[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  frequencyTotals_143 = _RAND_145[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  frequencyTotals_144 = _RAND_146[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  frequencyTotals_145 = _RAND_147[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  frequencyTotals_146 = _RAND_148[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  frequencyTotals_147 = _RAND_149[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  frequencyTotals_148 = _RAND_150[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  frequencyTotals_149 = _RAND_151[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  frequencyTotals_150 = _RAND_152[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  frequencyTotals_151 = _RAND_153[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  frequencyTotals_152 = _RAND_154[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  frequencyTotals_153 = _RAND_155[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  frequencyTotals_154 = _RAND_156[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  frequencyTotals_155 = _RAND_157[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  frequencyTotals_156 = _RAND_158[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  frequencyTotals_157 = _RAND_159[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  frequencyTotals_158 = _RAND_160[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  frequencyTotals_159 = _RAND_161[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  frequencyTotals_160 = _RAND_162[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  frequencyTotals_161 = _RAND_163[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  frequencyTotals_162 = _RAND_164[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  frequencyTotals_163 = _RAND_165[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  frequencyTotals_164 = _RAND_166[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  frequencyTotals_165 = _RAND_167[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  frequencyTotals_166 = _RAND_168[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  frequencyTotals_167 = _RAND_169[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  frequencyTotals_168 = _RAND_170[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  frequencyTotals_169 = _RAND_171[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  frequencyTotals_170 = _RAND_172[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  frequencyTotals_171 = _RAND_173[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  frequencyTotals_172 = _RAND_174[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  frequencyTotals_173 = _RAND_175[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  frequencyTotals_174 = _RAND_176[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  frequencyTotals_175 = _RAND_177[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  frequencyTotals_176 = _RAND_178[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  frequencyTotals_177 = _RAND_179[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  frequencyTotals_178 = _RAND_180[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  frequencyTotals_179 = _RAND_181[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  frequencyTotals_180 = _RAND_182[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  frequencyTotals_181 = _RAND_183[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  frequencyTotals_182 = _RAND_184[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  frequencyTotals_183 = _RAND_185[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  frequencyTotals_184 = _RAND_186[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  frequencyTotals_185 = _RAND_187[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  frequencyTotals_186 = _RAND_188[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  frequencyTotals_187 = _RAND_189[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  frequencyTotals_188 = _RAND_190[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  frequencyTotals_189 = _RAND_191[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  frequencyTotals_190 = _RAND_192[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  frequencyTotals_191 = _RAND_193[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  frequencyTotals_192 = _RAND_194[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  frequencyTotals_193 = _RAND_195[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  frequencyTotals_194 = _RAND_196[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  frequencyTotals_195 = _RAND_197[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  frequencyTotals_196 = _RAND_198[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  frequencyTotals_197 = _RAND_199[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  frequencyTotals_198 = _RAND_200[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  frequencyTotals_199 = _RAND_201[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  frequencyTotals_200 = _RAND_202[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  frequencyTotals_201 = _RAND_203[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  frequencyTotals_202 = _RAND_204[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  frequencyTotals_203 = _RAND_205[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  frequencyTotals_204 = _RAND_206[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  frequencyTotals_205 = _RAND_207[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  frequencyTotals_206 = _RAND_208[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  frequencyTotals_207 = _RAND_209[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  frequencyTotals_208 = _RAND_210[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  frequencyTotals_209 = _RAND_211[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  frequencyTotals_210 = _RAND_212[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  frequencyTotals_211 = _RAND_213[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  frequencyTotals_212 = _RAND_214[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  frequencyTotals_213 = _RAND_215[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  frequencyTotals_214 = _RAND_216[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  frequencyTotals_215 = _RAND_217[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  frequencyTotals_216 = _RAND_218[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  frequencyTotals_217 = _RAND_219[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  frequencyTotals_218 = _RAND_220[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  frequencyTotals_219 = _RAND_221[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  frequencyTotals_220 = _RAND_222[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  frequencyTotals_221 = _RAND_223[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  frequencyTotals_222 = _RAND_224[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  frequencyTotals_223 = _RAND_225[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  frequencyTotals_224 = _RAND_226[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  frequencyTotals_225 = _RAND_227[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  frequencyTotals_226 = _RAND_228[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  frequencyTotals_227 = _RAND_229[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  frequencyTotals_228 = _RAND_230[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  frequencyTotals_229 = _RAND_231[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  frequencyTotals_230 = _RAND_232[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  frequencyTotals_231 = _RAND_233[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  frequencyTotals_232 = _RAND_234[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  frequencyTotals_233 = _RAND_235[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  frequencyTotals_234 = _RAND_236[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  frequencyTotals_235 = _RAND_237[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  frequencyTotals_236 = _RAND_238[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  frequencyTotals_237 = _RAND_239[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  frequencyTotals_238 = _RAND_240[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  frequencyTotals_239 = _RAND_241[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  frequencyTotals_240 = _RAND_242[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  frequencyTotals_241 = _RAND_243[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  frequencyTotals_242 = _RAND_244[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  frequencyTotals_243 = _RAND_245[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  frequencyTotals_244 = _RAND_246[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  frequencyTotals_245 = _RAND_247[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  frequencyTotals_246 = _RAND_248[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  frequencyTotals_247 = _RAND_249[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  frequencyTotals_248 = _RAND_250[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  frequencyTotals_249 = _RAND_251[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  frequencyTotals_250 = _RAND_252[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  frequencyTotals_251 = _RAND_253[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  frequencyTotals_252 = _RAND_254[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  frequencyTotals_253 = _RAND_255[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  frequencyTotals_254 = _RAND_256[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  frequencyTotals_255 = _RAND_257[12:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else if (_T) begin
      state <= _GEN_1;
    end else if (state) begin
      if (io_dataIn_ready) begin
        if (_T_773) begin
          state <= 1'h0;
        end
      end
    end
    if (_T) begin
      if (io_start) begin
        currentByte <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        currentByte <= _T_772;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_0 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_0 <= _T_5;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_1 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_1 <= _T_8;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_2 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_2 <= _T_11;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_3 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_3 <= _T_14;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_4 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_4 <= _T_17;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_5 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_5 <= _T_20;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_6 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_6 <= _T_23;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_7 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_7 <= _T_26;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_8 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_8 <= _T_29;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_9 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_9 <= _T_32;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_10 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_10 <= _T_35;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_11 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_11 <= _T_38;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_12 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_12 <= _T_41;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_13 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_13 <= _T_44;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_14 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_14 <= _T_47;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_15 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_15 <= _T_50;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_16 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_16 <= _T_53;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_17 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_17 <= _T_56;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_18 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_18 <= _T_59;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_19 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_19 <= _T_62;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_20 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_20 <= _T_65;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_21 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_21 <= _T_68;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_22 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_22 <= _T_71;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_23 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_23 <= _T_74;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_24 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_24 <= _T_77;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_25 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_25 <= _T_80;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_26 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_26 <= _T_83;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_27 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_27 <= _T_86;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_28 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_28 <= _T_89;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_29 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_29 <= _T_92;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_30 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_30 <= _T_95;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_31 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_31 <= _T_98;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_32 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_32 <= _T_101;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_33 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_33 <= _T_104;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_34 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_34 <= _T_107;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_35 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_35 <= _T_110;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_36 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_36 <= _T_113;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_37 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_37 <= _T_116;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_38 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_38 <= _T_119;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_39 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_39 <= _T_122;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_40 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_40 <= _T_125;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_41 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_41 <= _T_128;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_42 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_42 <= _T_131;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_43 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_43 <= _T_134;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_44 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_44 <= _T_137;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_45 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_45 <= _T_140;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_46 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_46 <= _T_143;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_47 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_47 <= _T_146;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_48 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_48 <= _T_149;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_49 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_49 <= _T_152;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_50 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_50 <= _T_155;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_51 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_51 <= _T_158;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_52 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_52 <= _T_161;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_53 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_53 <= _T_164;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_54 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_54 <= _T_167;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_55 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_55 <= _T_170;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_56 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_56 <= _T_173;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_57 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_57 <= _T_176;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_58 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_58 <= _T_179;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_59 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_59 <= _T_182;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_60 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_60 <= _T_185;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_61 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_61 <= _T_188;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_62 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_62 <= _T_191;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_63 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_63 <= _T_194;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_64 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_64 <= _T_197;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_65 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_65 <= _T_200;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_66 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_66 <= _T_203;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_67 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_67 <= _T_206;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_68 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_68 <= _T_209;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_69 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_69 <= _T_212;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_70 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_70 <= _T_215;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_71 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_71 <= _T_218;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_72 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_72 <= _T_221;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_73 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_73 <= _T_224;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_74 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_74 <= _T_227;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_75 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_75 <= _T_230;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_76 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_76 <= _T_233;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_77 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_77 <= _T_236;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_78 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_78 <= _T_239;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_79 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_79 <= _T_242;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_80 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_80 <= _T_245;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_81 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_81 <= _T_248;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_82 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_82 <= _T_251;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_83 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_83 <= _T_254;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_84 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_84 <= _T_257;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_85 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_85 <= _T_260;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_86 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_86 <= _T_263;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_87 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_87 <= _T_266;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_88 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_88 <= _T_269;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_89 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_89 <= _T_272;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_90 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_90 <= _T_275;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_91 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_91 <= _T_278;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_92 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_92 <= _T_281;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_93 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_93 <= _T_284;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_94 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_94 <= _T_287;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_95 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_95 <= _T_290;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_96 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_96 <= _T_293;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_97 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_97 <= _T_296;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_98 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_98 <= _T_299;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_99 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_99 <= _T_302;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_100 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_100 <= _T_305;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_101 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_101 <= _T_308;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_102 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_102 <= _T_311;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_103 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_103 <= _T_314;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_104 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_104 <= _T_317;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_105 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_105 <= _T_320;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_106 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_106 <= _T_323;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_107 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_107 <= _T_326;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_108 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_108 <= _T_329;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_109 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_109 <= _T_332;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_110 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_110 <= _T_335;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_111 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_111 <= _T_338;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_112 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_112 <= _T_341;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_113 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_113 <= _T_344;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_114 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_114 <= _T_347;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_115 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_115 <= _T_350;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_116 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_116 <= _T_353;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_117 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_117 <= _T_356;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_118 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_118 <= _T_359;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_119 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_119 <= _T_362;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_120 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_120 <= _T_365;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_121 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_121 <= _T_368;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_122 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_122 <= _T_371;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_123 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_123 <= _T_374;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_124 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_124 <= _T_377;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_125 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_125 <= _T_380;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_126 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_126 <= _T_383;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_127 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_127 <= _T_386;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_128 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_128 <= _T_389;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_129 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_129 <= _T_392;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_130 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_130 <= _T_395;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_131 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_131 <= _T_398;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_132 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_132 <= _T_401;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_133 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_133 <= _T_404;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_134 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_134 <= _T_407;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_135 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_135 <= _T_410;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_136 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_136 <= _T_413;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_137 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_137 <= _T_416;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_138 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_138 <= _T_419;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_139 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_139 <= _T_422;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_140 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_140 <= _T_425;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_141 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_141 <= _T_428;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_142 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_142 <= _T_431;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_143 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_143 <= _T_434;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_144 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_144 <= _T_437;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_145 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_145 <= _T_440;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_146 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_146 <= _T_443;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_147 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_147 <= _T_446;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_148 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_148 <= _T_449;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_149 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_149 <= _T_452;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_150 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_150 <= _T_455;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_151 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_151 <= _T_458;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_152 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_152 <= _T_461;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_153 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_153 <= _T_464;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_154 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_154 <= _T_467;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_155 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_155 <= _T_470;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_156 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_156 <= _T_473;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_157 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_157 <= _T_476;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_158 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_158 <= _T_479;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_159 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_159 <= _T_482;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_160 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_160 <= _T_485;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_161 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_161 <= _T_488;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_162 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_162 <= _T_491;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_163 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_163 <= _T_494;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_164 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_164 <= _T_497;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_165 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_165 <= _T_500;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_166 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_166 <= _T_503;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_167 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_167 <= _T_506;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_168 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_168 <= _T_509;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_169 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_169 <= _T_512;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_170 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_170 <= _T_515;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_171 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_171 <= _T_518;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_172 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_172 <= _T_521;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_173 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_173 <= _T_524;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_174 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_174 <= _T_527;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_175 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_175 <= _T_530;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_176 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_176 <= _T_533;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_177 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_177 <= _T_536;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_178 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_178 <= _T_539;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_179 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_179 <= _T_542;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_180 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_180 <= _T_545;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_181 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_181 <= _T_548;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_182 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_182 <= _T_551;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_183 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_183 <= _T_554;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_184 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_184 <= _T_557;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_185 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_185 <= _T_560;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_186 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_186 <= _T_563;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_187 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_187 <= _T_566;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_188 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_188 <= _T_569;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_189 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_189 <= _T_572;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_190 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_190 <= _T_575;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_191 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_191 <= _T_578;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_192 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_192 <= _T_581;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_193 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_193 <= _T_584;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_194 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_194 <= _T_587;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_195 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_195 <= _T_590;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_196 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_196 <= _T_593;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_197 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_197 <= _T_596;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_198 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_198 <= _T_599;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_199 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_199 <= _T_602;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_200 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_200 <= _T_605;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_201 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_201 <= _T_608;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_202 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_202 <= _T_611;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_203 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_203 <= _T_614;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_204 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_204 <= _T_617;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_205 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_205 <= _T_620;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_206 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_206 <= _T_623;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_207 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_207 <= _T_626;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_208 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_208 <= _T_629;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_209 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_209 <= _T_632;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_210 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_210 <= _T_635;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_211 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_211 <= _T_638;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_212 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_212 <= _T_641;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_213 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_213 <= _T_644;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_214 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_214 <= _T_647;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_215 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_215 <= _T_650;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_216 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_216 <= _T_653;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_217 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_217 <= _T_656;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_218 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_218 <= _T_659;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_219 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_219 <= _T_662;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_220 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_220 <= _T_665;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_221 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_221 <= _T_668;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_222 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_222 <= _T_671;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_223 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_223 <= _T_674;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_224 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_224 <= _T_677;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_225 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_225 <= _T_680;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_226 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_226 <= _T_683;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_227 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_227 <= _T_686;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_228 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_228 <= _T_689;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_229 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_229 <= _T_692;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_230 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_230 <= _T_695;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_231 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_231 <= _T_698;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_232 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_232 <= _T_701;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_233 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_233 <= _T_704;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_234 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_234 <= _T_707;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_235 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_235 <= _T_710;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_236 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_236 <= _T_713;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_237 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_237 <= _T_716;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_238 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_238 <= _T_719;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_239 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_239 <= _T_722;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_240 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_240 <= _T_725;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_241 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_241 <= _T_728;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_242 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_242 <= _T_731;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_243 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_243 <= _T_734;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_244 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_244 <= _T_737;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_245 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_245 <= _T_740;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_246 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_246 <= _T_743;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_247 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_247 <= _T_746;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_248 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_248 <= _T_749;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_249 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_249 <= _T_752;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_250 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_250 <= _T_755;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_251 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_251 <= _T_758;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_252 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_252 <= _T_761;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_253 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_253 <= _T_764;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_254 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_254 <= _T_767;
      end
    end
    if (_T) begin
      if (io_start) begin
        frequencyTotals_255 <= 13'h0;
      end
    end else if (state) begin
      if (io_dataIn_ready) begin
        frequencyTotals_255 <= _T_770;
      end
    end
  end
endmodule
module characterFrequencySort(
  input         clock,
  input         reset,
  input         io_start,
  input  [12:0] io_dataIn_0,
  input  [12:0] io_dataIn_1,
  input  [12:0] io_dataIn_2,
  input  [12:0] io_dataIn_3,
  input  [12:0] io_dataIn_4,
  input  [12:0] io_dataIn_5,
  input  [12:0] io_dataIn_6,
  input  [12:0] io_dataIn_7,
  input  [12:0] io_dataIn_8,
  input  [12:0] io_dataIn_9,
  input  [12:0] io_dataIn_10,
  input  [12:0] io_dataIn_11,
  input  [12:0] io_dataIn_12,
  input  [12:0] io_dataIn_13,
  input  [12:0] io_dataIn_14,
  input  [12:0] io_dataIn_15,
  input  [12:0] io_dataIn_16,
  input  [12:0] io_dataIn_17,
  input  [12:0] io_dataIn_18,
  input  [12:0] io_dataIn_19,
  input  [12:0] io_dataIn_20,
  input  [12:0] io_dataIn_21,
  input  [12:0] io_dataIn_22,
  input  [12:0] io_dataIn_23,
  input  [12:0] io_dataIn_24,
  input  [12:0] io_dataIn_25,
  input  [12:0] io_dataIn_26,
  input  [12:0] io_dataIn_27,
  input  [12:0] io_dataIn_28,
  input  [12:0] io_dataIn_29,
  input  [12:0] io_dataIn_30,
  input  [12:0] io_dataIn_31,
  input  [12:0] io_dataIn_32,
  input  [12:0] io_dataIn_33,
  input  [12:0] io_dataIn_34,
  input  [12:0] io_dataIn_35,
  input  [12:0] io_dataIn_36,
  input  [12:0] io_dataIn_37,
  input  [12:0] io_dataIn_38,
  input  [12:0] io_dataIn_39,
  input  [12:0] io_dataIn_40,
  input  [12:0] io_dataIn_41,
  input  [12:0] io_dataIn_42,
  input  [12:0] io_dataIn_43,
  input  [12:0] io_dataIn_44,
  input  [12:0] io_dataIn_45,
  input  [12:0] io_dataIn_46,
  input  [12:0] io_dataIn_47,
  input  [12:0] io_dataIn_48,
  input  [12:0] io_dataIn_49,
  input  [12:0] io_dataIn_50,
  input  [12:0] io_dataIn_51,
  input  [12:0] io_dataIn_52,
  input  [12:0] io_dataIn_53,
  input  [12:0] io_dataIn_54,
  input  [12:0] io_dataIn_55,
  input  [12:0] io_dataIn_56,
  input  [12:0] io_dataIn_57,
  input  [12:0] io_dataIn_58,
  input  [12:0] io_dataIn_59,
  input  [12:0] io_dataIn_60,
  input  [12:0] io_dataIn_61,
  input  [12:0] io_dataIn_62,
  input  [12:0] io_dataIn_63,
  input  [12:0] io_dataIn_64,
  input  [12:0] io_dataIn_65,
  input  [12:0] io_dataIn_66,
  input  [12:0] io_dataIn_67,
  input  [12:0] io_dataIn_68,
  input  [12:0] io_dataIn_69,
  input  [12:0] io_dataIn_70,
  input  [12:0] io_dataIn_71,
  input  [12:0] io_dataIn_72,
  input  [12:0] io_dataIn_73,
  input  [12:0] io_dataIn_74,
  input  [12:0] io_dataIn_75,
  input  [12:0] io_dataIn_76,
  input  [12:0] io_dataIn_77,
  input  [12:0] io_dataIn_78,
  input  [12:0] io_dataIn_79,
  input  [12:0] io_dataIn_80,
  input  [12:0] io_dataIn_81,
  input  [12:0] io_dataIn_82,
  input  [12:0] io_dataIn_83,
  input  [12:0] io_dataIn_84,
  input  [12:0] io_dataIn_85,
  input  [12:0] io_dataIn_86,
  input  [12:0] io_dataIn_87,
  input  [12:0] io_dataIn_88,
  input  [12:0] io_dataIn_89,
  input  [12:0] io_dataIn_90,
  input  [12:0] io_dataIn_91,
  input  [12:0] io_dataIn_92,
  input  [12:0] io_dataIn_93,
  input  [12:0] io_dataIn_94,
  input  [12:0] io_dataIn_95,
  input  [12:0] io_dataIn_96,
  input  [12:0] io_dataIn_97,
  input  [12:0] io_dataIn_98,
  input  [12:0] io_dataIn_99,
  input  [12:0] io_dataIn_100,
  input  [12:0] io_dataIn_101,
  input  [12:0] io_dataIn_102,
  input  [12:0] io_dataIn_103,
  input  [12:0] io_dataIn_104,
  input  [12:0] io_dataIn_105,
  input  [12:0] io_dataIn_106,
  input  [12:0] io_dataIn_107,
  input  [12:0] io_dataIn_108,
  input  [12:0] io_dataIn_109,
  input  [12:0] io_dataIn_110,
  input  [12:0] io_dataIn_111,
  input  [12:0] io_dataIn_112,
  input  [12:0] io_dataIn_113,
  input  [12:0] io_dataIn_114,
  input  [12:0] io_dataIn_115,
  input  [12:0] io_dataIn_116,
  input  [12:0] io_dataIn_117,
  input  [12:0] io_dataIn_118,
  input  [12:0] io_dataIn_119,
  input  [12:0] io_dataIn_120,
  input  [12:0] io_dataIn_121,
  input  [12:0] io_dataIn_122,
  input  [12:0] io_dataIn_123,
  input  [12:0] io_dataIn_124,
  input  [12:0] io_dataIn_125,
  input  [12:0] io_dataIn_126,
  input  [12:0] io_dataIn_127,
  input  [12:0] io_dataIn_128,
  input  [12:0] io_dataIn_129,
  input  [12:0] io_dataIn_130,
  input  [12:0] io_dataIn_131,
  input  [12:0] io_dataIn_132,
  input  [12:0] io_dataIn_133,
  input  [12:0] io_dataIn_134,
  input  [12:0] io_dataIn_135,
  input  [12:0] io_dataIn_136,
  input  [12:0] io_dataIn_137,
  input  [12:0] io_dataIn_138,
  input  [12:0] io_dataIn_139,
  input  [12:0] io_dataIn_140,
  input  [12:0] io_dataIn_141,
  input  [12:0] io_dataIn_142,
  input  [12:0] io_dataIn_143,
  input  [12:0] io_dataIn_144,
  input  [12:0] io_dataIn_145,
  input  [12:0] io_dataIn_146,
  input  [12:0] io_dataIn_147,
  input  [12:0] io_dataIn_148,
  input  [12:0] io_dataIn_149,
  input  [12:0] io_dataIn_150,
  input  [12:0] io_dataIn_151,
  input  [12:0] io_dataIn_152,
  input  [12:0] io_dataIn_153,
  input  [12:0] io_dataIn_154,
  input  [12:0] io_dataIn_155,
  input  [12:0] io_dataIn_156,
  input  [12:0] io_dataIn_157,
  input  [12:0] io_dataIn_158,
  input  [12:0] io_dataIn_159,
  input  [12:0] io_dataIn_160,
  input  [12:0] io_dataIn_161,
  input  [12:0] io_dataIn_162,
  input  [12:0] io_dataIn_163,
  input  [12:0] io_dataIn_164,
  input  [12:0] io_dataIn_165,
  input  [12:0] io_dataIn_166,
  input  [12:0] io_dataIn_167,
  input  [12:0] io_dataIn_168,
  input  [12:0] io_dataIn_169,
  input  [12:0] io_dataIn_170,
  input  [12:0] io_dataIn_171,
  input  [12:0] io_dataIn_172,
  input  [12:0] io_dataIn_173,
  input  [12:0] io_dataIn_174,
  input  [12:0] io_dataIn_175,
  input  [12:0] io_dataIn_176,
  input  [12:0] io_dataIn_177,
  input  [12:0] io_dataIn_178,
  input  [12:0] io_dataIn_179,
  input  [12:0] io_dataIn_180,
  input  [12:0] io_dataIn_181,
  input  [12:0] io_dataIn_182,
  input  [12:0] io_dataIn_183,
  input  [12:0] io_dataIn_184,
  input  [12:0] io_dataIn_185,
  input  [12:0] io_dataIn_186,
  input  [12:0] io_dataIn_187,
  input  [12:0] io_dataIn_188,
  input  [12:0] io_dataIn_189,
  input  [12:0] io_dataIn_190,
  input  [12:0] io_dataIn_191,
  input  [12:0] io_dataIn_192,
  input  [12:0] io_dataIn_193,
  input  [12:0] io_dataIn_194,
  input  [12:0] io_dataIn_195,
  input  [12:0] io_dataIn_196,
  input  [12:0] io_dataIn_197,
  input  [12:0] io_dataIn_198,
  input  [12:0] io_dataIn_199,
  input  [12:0] io_dataIn_200,
  input  [12:0] io_dataIn_201,
  input  [12:0] io_dataIn_202,
  input  [12:0] io_dataIn_203,
  input  [12:0] io_dataIn_204,
  input  [12:0] io_dataIn_205,
  input  [12:0] io_dataIn_206,
  input  [12:0] io_dataIn_207,
  input  [12:0] io_dataIn_208,
  input  [12:0] io_dataIn_209,
  input  [12:0] io_dataIn_210,
  input  [12:0] io_dataIn_211,
  input  [12:0] io_dataIn_212,
  input  [12:0] io_dataIn_213,
  input  [12:0] io_dataIn_214,
  input  [12:0] io_dataIn_215,
  input  [12:0] io_dataIn_216,
  input  [12:0] io_dataIn_217,
  input  [12:0] io_dataIn_218,
  input  [12:0] io_dataIn_219,
  input  [12:0] io_dataIn_220,
  input  [12:0] io_dataIn_221,
  input  [12:0] io_dataIn_222,
  input  [12:0] io_dataIn_223,
  input  [12:0] io_dataIn_224,
  input  [12:0] io_dataIn_225,
  input  [12:0] io_dataIn_226,
  input  [12:0] io_dataIn_227,
  input  [12:0] io_dataIn_228,
  input  [12:0] io_dataIn_229,
  input  [12:0] io_dataIn_230,
  input  [12:0] io_dataIn_231,
  input  [12:0] io_dataIn_232,
  input  [12:0] io_dataIn_233,
  input  [12:0] io_dataIn_234,
  input  [12:0] io_dataIn_235,
  input  [12:0] io_dataIn_236,
  input  [12:0] io_dataIn_237,
  input  [12:0] io_dataIn_238,
  input  [12:0] io_dataIn_239,
  input  [12:0] io_dataIn_240,
  input  [12:0] io_dataIn_241,
  input  [12:0] io_dataIn_242,
  input  [12:0] io_dataIn_243,
  input  [12:0] io_dataIn_244,
  input  [12:0] io_dataIn_245,
  input  [12:0] io_dataIn_246,
  input  [12:0] io_dataIn_247,
  input  [12:0] io_dataIn_248,
  input  [12:0] io_dataIn_249,
  input  [12:0] io_dataIn_250,
  input  [12:0] io_dataIn_251,
  input  [12:0] io_dataIn_252,
  input  [12:0] io_dataIn_253,
  input  [12:0] io_dataIn_254,
  input  [12:0] io_dataIn_255,
  output [12:0] io_sortedFrequency_0,
  output [12:0] io_sortedFrequency_1,
  output [12:0] io_sortedFrequency_2,
  output [12:0] io_sortedFrequency_3,
  output [12:0] io_sortedFrequency_4,
  output [12:0] io_sortedFrequency_5,
  output [12:0] io_sortedFrequency_6,
  output [12:0] io_sortedFrequency_7,
  output [12:0] io_sortedFrequency_8,
  output [12:0] io_sortedFrequency_9,
  output [12:0] io_sortedFrequency_10,
  output [12:0] io_sortedFrequency_11,
  output [12:0] io_sortedFrequency_12,
  output [12:0] io_sortedFrequency_13,
  output [12:0] io_sortedFrequency_14,
  output [12:0] io_sortedFrequency_15,
  output [12:0] io_sortedFrequency_16,
  output [12:0] io_sortedFrequency_17,
  output [12:0] io_sortedFrequency_18,
  output [12:0] io_sortedFrequency_19,
  output [12:0] io_sortedFrequency_20,
  output [12:0] io_sortedFrequency_21,
  output [12:0] io_sortedFrequency_22,
  output [12:0] io_sortedFrequency_23,
  output [12:0] io_sortedFrequency_24,
  output [12:0] io_sortedFrequency_25,
  output [12:0] io_sortedFrequency_26,
  output [12:0] io_sortedFrequency_27,
  output [12:0] io_sortedFrequency_28,
  output [12:0] io_sortedFrequency_29,
  output [12:0] io_sortedFrequency_30,
  output [12:0] io_sortedFrequency_31,
  output [8:0]  io_sortedCharacter_0,
  output [8:0]  io_sortedCharacter_1,
  output [8:0]  io_sortedCharacter_2,
  output [8:0]  io_sortedCharacter_3,
  output [8:0]  io_sortedCharacter_4,
  output [8:0]  io_sortedCharacter_5,
  output [8:0]  io_sortedCharacter_6,
  output [8:0]  io_sortedCharacter_7,
  output [8:0]  io_sortedCharacter_8,
  output [8:0]  io_sortedCharacter_9,
  output [8:0]  io_sortedCharacter_10,
  output [8:0]  io_sortedCharacter_11,
  output [8:0]  io_sortedCharacter_12,
  output [8:0]  io_sortedCharacter_13,
  output [8:0]  io_sortedCharacter_14,
  output [8:0]  io_sortedCharacter_15,
  output [8:0]  io_sortedCharacter_16,
  output [8:0]  io_sortedCharacter_17,
  output [8:0]  io_sortedCharacter_18,
  output [8:0]  io_sortedCharacter_19,
  output [8:0]  io_sortedCharacter_20,
  output [8:0]  io_sortedCharacter_21,
  output [8:0]  io_sortedCharacter_22,
  output [8:0]  io_sortedCharacter_23,
  output [8:0]  io_sortedCharacter_24,
  output [8:0]  io_sortedCharacter_25,
  output [8:0]  io_sortedCharacter_26,
  output [8:0]  io_sortedCharacter_27,
  output [8:0]  io_sortedCharacter_28,
  output [8:0]  io_sortedCharacter_29,
  output [8:0]  io_sortedCharacter_30,
  output [8:0]  io_sortedCharacter_31,
  output        io_finished
);
  reg [1:0] state; // @[characterFrequencySort.scala 23:22]
  reg [31:0] _RAND_0;
  reg [8:0] iteration; // @[characterFrequencySort.scala 31:22]
  reg [31:0] _RAND_1;
  reg [12:0] sortedFrequency_0; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_2;
  reg [12:0] sortedFrequency_1; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_3;
  reg [12:0] sortedFrequency_2; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_4;
  reg [12:0] sortedFrequency_3; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_5;
  reg [12:0] sortedFrequency_4; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_6;
  reg [12:0] sortedFrequency_5; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_7;
  reg [12:0] sortedFrequency_6; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_8;
  reg [12:0] sortedFrequency_7; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_9;
  reg [12:0] sortedFrequency_8; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_10;
  reg [12:0] sortedFrequency_9; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_11;
  reg [12:0] sortedFrequency_10; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_12;
  reg [12:0] sortedFrequency_11; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_13;
  reg [12:0] sortedFrequency_12; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_14;
  reg [12:0] sortedFrequency_13; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_15;
  reg [12:0] sortedFrequency_14; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_16;
  reg [12:0] sortedFrequency_15; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_17;
  reg [12:0] sortedFrequency_16; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_18;
  reg [12:0] sortedFrequency_17; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_19;
  reg [12:0] sortedFrequency_18; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_20;
  reg [12:0] sortedFrequency_19; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_21;
  reg [12:0] sortedFrequency_20; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_22;
  reg [12:0] sortedFrequency_21; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_23;
  reg [12:0] sortedFrequency_22; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_24;
  reg [12:0] sortedFrequency_23; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_25;
  reg [12:0] sortedFrequency_24; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_26;
  reg [12:0] sortedFrequency_25; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_27;
  reg [12:0] sortedFrequency_26; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_28;
  reg [12:0] sortedFrequency_27; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_29;
  reg [12:0] sortedFrequency_28; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_30;
  reg [12:0] sortedFrequency_29; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_31;
  reg [12:0] sortedFrequency_30; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_32;
  reg [12:0] sortedFrequency_31; // @[characterFrequencySort.scala 34:28]
  reg [31:0] _RAND_33;
  reg [8:0] sortedCharacter_0; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_34;
  reg [8:0] sortedCharacter_1; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_35;
  reg [8:0] sortedCharacter_2; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_36;
  reg [8:0] sortedCharacter_3; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_37;
  reg [8:0] sortedCharacter_4; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_38;
  reg [8:0] sortedCharacter_5; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_39;
  reg [8:0] sortedCharacter_6; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_40;
  reg [8:0] sortedCharacter_7; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_41;
  reg [8:0] sortedCharacter_8; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_42;
  reg [8:0] sortedCharacter_9; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_43;
  reg [8:0] sortedCharacter_10; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_44;
  reg [8:0] sortedCharacter_11; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_45;
  reg [8:0] sortedCharacter_12; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_46;
  reg [8:0] sortedCharacter_13; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_47;
  reg [8:0] sortedCharacter_14; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_48;
  reg [8:0] sortedCharacter_15; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_49;
  reg [8:0] sortedCharacter_16; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_50;
  reg [8:0] sortedCharacter_17; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_51;
  reg [8:0] sortedCharacter_18; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_52;
  reg [8:0] sortedCharacter_19; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_53;
  reg [8:0] sortedCharacter_20; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_54;
  reg [8:0] sortedCharacter_21; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_55;
  reg [8:0] sortedCharacter_22; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_56;
  reg [8:0] sortedCharacter_23; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_57;
  reg [8:0] sortedCharacter_24; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_58;
  reg [8:0] sortedCharacter_25; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_59;
  reg [8:0] sortedCharacter_26; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_60;
  reg [8:0] sortedCharacter_27; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_61;
  reg [8:0] sortedCharacter_28; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_62;
  reg [8:0] sortedCharacter_29; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_63;
  reg [8:0] sortedCharacter_30; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_64;
  reg [8:0] sortedCharacter_31; // @[characterFrequencySort.scala 35:28]
  reg [31:0] _RAND_65;
  reg [12:0] sortedFrequencyTemp_0; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_66;
  reg [12:0] sortedFrequencyTemp_1; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_67;
  reg [12:0] sortedFrequencyTemp_2; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_68;
  reg [12:0] sortedFrequencyTemp_3; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_69;
  reg [12:0] sortedFrequencyTemp_4; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_70;
  reg [12:0] sortedFrequencyTemp_5; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_71;
  reg [12:0] sortedFrequencyTemp_6; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_72;
  reg [12:0] sortedFrequencyTemp_7; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_73;
  reg [12:0] sortedFrequencyTemp_8; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_74;
  reg [12:0] sortedFrequencyTemp_9; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_75;
  reg [12:0] sortedFrequencyTemp_10; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_76;
  reg [12:0] sortedFrequencyTemp_11; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_77;
  reg [12:0] sortedFrequencyTemp_12; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_78;
  reg [12:0] sortedFrequencyTemp_13; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_79;
  reg [12:0] sortedFrequencyTemp_14; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_80;
  reg [12:0] sortedFrequencyTemp_15; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_81;
  reg [12:0] sortedFrequencyTemp_16; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_82;
  reg [12:0] sortedFrequencyTemp_17; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_83;
  reg [12:0] sortedFrequencyTemp_18; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_84;
  reg [12:0] sortedFrequencyTemp_19; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_85;
  reg [12:0] sortedFrequencyTemp_20; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_86;
  reg [12:0] sortedFrequencyTemp_21; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_87;
  reg [12:0] sortedFrequencyTemp_22; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_88;
  reg [12:0] sortedFrequencyTemp_23; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_89;
  reg [12:0] sortedFrequencyTemp_24; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_90;
  reg [12:0] sortedFrequencyTemp_25; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_91;
  reg [12:0] sortedFrequencyTemp_26; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_92;
  reg [12:0] sortedFrequencyTemp_27; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_93;
  reg [12:0] sortedFrequencyTemp_28; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_94;
  reg [12:0] sortedFrequencyTemp_29; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_95;
  reg [12:0] sortedFrequencyTemp_30; // @[characterFrequencySort.scala 37:32]
  reg [31:0] _RAND_96;
  reg [8:0] sortedCharacterTemp_0; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_97;
  reg [8:0] sortedCharacterTemp_1; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_98;
  reg [8:0] sortedCharacterTemp_2; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_99;
  reg [8:0] sortedCharacterTemp_3; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_100;
  reg [8:0] sortedCharacterTemp_4; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_101;
  reg [8:0] sortedCharacterTemp_5; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_102;
  reg [8:0] sortedCharacterTemp_6; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_103;
  reg [8:0] sortedCharacterTemp_7; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_104;
  reg [8:0] sortedCharacterTemp_8; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_105;
  reg [8:0] sortedCharacterTemp_9; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_106;
  reg [8:0] sortedCharacterTemp_10; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_107;
  reg [8:0] sortedCharacterTemp_11; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_108;
  reg [8:0] sortedCharacterTemp_12; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_109;
  reg [8:0] sortedCharacterTemp_13; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_110;
  reg [8:0] sortedCharacterTemp_14; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_111;
  reg [8:0] sortedCharacterTemp_15; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_112;
  reg [8:0] sortedCharacterTemp_16; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_113;
  reg [8:0] sortedCharacterTemp_17; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_114;
  reg [8:0] sortedCharacterTemp_18; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_115;
  reg [8:0] sortedCharacterTemp_19; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_116;
  reg [8:0] sortedCharacterTemp_20; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_117;
  reg [8:0] sortedCharacterTemp_21; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_118;
  reg [8:0] sortedCharacterTemp_22; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_119;
  reg [8:0] sortedCharacterTemp_23; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_120;
  reg [8:0] sortedCharacterTemp_24; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_121;
  reg [8:0] sortedCharacterTemp_25; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_122;
  reg [8:0] sortedCharacterTemp_26; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_123;
  reg [8:0] sortedCharacterTemp_27; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_124;
  reg [8:0] sortedCharacterTemp_28; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_125;
  reg [8:0] sortedCharacterTemp_29; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_126;
  reg [8:0] sortedCharacterTemp_30; // @[characterFrequencySort.scala 38:32]
  reg [31:0] _RAND_127;
  reg [12:0] escapeFrequency; // @[characterFrequencySort.scala 42:28]
  reg [31:0] _RAND_128;
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire [15:0] _GEN_987 = {{7'd0}, iteration}; // @[characterFrequencySort.scala 66:22]
  wire  _T_6 = _GEN_987 < 16'h100; // @[characterFrequencySort.scala 66:22]
  wire [12:0] _GEN_68 = 8'h1 == iteration[7:0] ? io_dataIn_1 : io_dataIn_0; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_69 = 8'h2 == iteration[7:0] ? io_dataIn_2 : _GEN_68; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_70 = 8'h3 == iteration[7:0] ? io_dataIn_3 : _GEN_69; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_71 = 8'h4 == iteration[7:0] ? io_dataIn_4 : _GEN_70; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_72 = 8'h5 == iteration[7:0] ? io_dataIn_5 : _GEN_71; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_73 = 8'h6 == iteration[7:0] ? io_dataIn_6 : _GEN_72; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_74 = 8'h7 == iteration[7:0] ? io_dataIn_7 : _GEN_73; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_75 = 8'h8 == iteration[7:0] ? io_dataIn_8 : _GEN_74; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_76 = 8'h9 == iteration[7:0] ? io_dataIn_9 : _GEN_75; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_77 = 8'ha == iteration[7:0] ? io_dataIn_10 : _GEN_76; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_78 = 8'hb == iteration[7:0] ? io_dataIn_11 : _GEN_77; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_79 = 8'hc == iteration[7:0] ? io_dataIn_12 : _GEN_78; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_80 = 8'hd == iteration[7:0] ? io_dataIn_13 : _GEN_79; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_81 = 8'he == iteration[7:0] ? io_dataIn_14 : _GEN_80; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_82 = 8'hf == iteration[7:0] ? io_dataIn_15 : _GEN_81; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_83 = 8'h10 == iteration[7:0] ? io_dataIn_16 : _GEN_82; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_84 = 8'h11 == iteration[7:0] ? io_dataIn_17 : _GEN_83; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_85 = 8'h12 == iteration[7:0] ? io_dataIn_18 : _GEN_84; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_86 = 8'h13 == iteration[7:0] ? io_dataIn_19 : _GEN_85; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_87 = 8'h14 == iteration[7:0] ? io_dataIn_20 : _GEN_86; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_88 = 8'h15 == iteration[7:0] ? io_dataIn_21 : _GEN_87; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_89 = 8'h16 == iteration[7:0] ? io_dataIn_22 : _GEN_88; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_90 = 8'h17 == iteration[7:0] ? io_dataIn_23 : _GEN_89; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_91 = 8'h18 == iteration[7:0] ? io_dataIn_24 : _GEN_90; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_92 = 8'h19 == iteration[7:0] ? io_dataIn_25 : _GEN_91; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_93 = 8'h1a == iteration[7:0] ? io_dataIn_26 : _GEN_92; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_94 = 8'h1b == iteration[7:0] ? io_dataIn_27 : _GEN_93; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_95 = 8'h1c == iteration[7:0] ? io_dataIn_28 : _GEN_94; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_96 = 8'h1d == iteration[7:0] ? io_dataIn_29 : _GEN_95; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_97 = 8'h1e == iteration[7:0] ? io_dataIn_30 : _GEN_96; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_98 = 8'h1f == iteration[7:0] ? io_dataIn_31 : _GEN_97; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_99 = 8'h20 == iteration[7:0] ? io_dataIn_32 : _GEN_98; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_100 = 8'h21 == iteration[7:0] ? io_dataIn_33 : _GEN_99; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_101 = 8'h22 == iteration[7:0] ? io_dataIn_34 : _GEN_100; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_102 = 8'h23 == iteration[7:0] ? io_dataIn_35 : _GEN_101; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_103 = 8'h24 == iteration[7:0] ? io_dataIn_36 : _GEN_102; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_104 = 8'h25 == iteration[7:0] ? io_dataIn_37 : _GEN_103; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_105 = 8'h26 == iteration[7:0] ? io_dataIn_38 : _GEN_104; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_106 = 8'h27 == iteration[7:0] ? io_dataIn_39 : _GEN_105; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_107 = 8'h28 == iteration[7:0] ? io_dataIn_40 : _GEN_106; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_108 = 8'h29 == iteration[7:0] ? io_dataIn_41 : _GEN_107; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_109 = 8'h2a == iteration[7:0] ? io_dataIn_42 : _GEN_108; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_110 = 8'h2b == iteration[7:0] ? io_dataIn_43 : _GEN_109; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_111 = 8'h2c == iteration[7:0] ? io_dataIn_44 : _GEN_110; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_112 = 8'h2d == iteration[7:0] ? io_dataIn_45 : _GEN_111; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_113 = 8'h2e == iteration[7:0] ? io_dataIn_46 : _GEN_112; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_114 = 8'h2f == iteration[7:0] ? io_dataIn_47 : _GEN_113; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_115 = 8'h30 == iteration[7:0] ? io_dataIn_48 : _GEN_114; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_116 = 8'h31 == iteration[7:0] ? io_dataIn_49 : _GEN_115; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_117 = 8'h32 == iteration[7:0] ? io_dataIn_50 : _GEN_116; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_118 = 8'h33 == iteration[7:0] ? io_dataIn_51 : _GEN_117; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_119 = 8'h34 == iteration[7:0] ? io_dataIn_52 : _GEN_118; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_120 = 8'h35 == iteration[7:0] ? io_dataIn_53 : _GEN_119; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_121 = 8'h36 == iteration[7:0] ? io_dataIn_54 : _GEN_120; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_122 = 8'h37 == iteration[7:0] ? io_dataIn_55 : _GEN_121; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_123 = 8'h38 == iteration[7:0] ? io_dataIn_56 : _GEN_122; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_124 = 8'h39 == iteration[7:0] ? io_dataIn_57 : _GEN_123; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_125 = 8'h3a == iteration[7:0] ? io_dataIn_58 : _GEN_124; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_126 = 8'h3b == iteration[7:0] ? io_dataIn_59 : _GEN_125; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_127 = 8'h3c == iteration[7:0] ? io_dataIn_60 : _GEN_126; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_128 = 8'h3d == iteration[7:0] ? io_dataIn_61 : _GEN_127; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_129 = 8'h3e == iteration[7:0] ? io_dataIn_62 : _GEN_128; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_130 = 8'h3f == iteration[7:0] ? io_dataIn_63 : _GEN_129; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_131 = 8'h40 == iteration[7:0] ? io_dataIn_64 : _GEN_130; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_132 = 8'h41 == iteration[7:0] ? io_dataIn_65 : _GEN_131; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_133 = 8'h42 == iteration[7:0] ? io_dataIn_66 : _GEN_132; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_134 = 8'h43 == iteration[7:0] ? io_dataIn_67 : _GEN_133; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_135 = 8'h44 == iteration[7:0] ? io_dataIn_68 : _GEN_134; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_136 = 8'h45 == iteration[7:0] ? io_dataIn_69 : _GEN_135; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_137 = 8'h46 == iteration[7:0] ? io_dataIn_70 : _GEN_136; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_138 = 8'h47 == iteration[7:0] ? io_dataIn_71 : _GEN_137; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_139 = 8'h48 == iteration[7:0] ? io_dataIn_72 : _GEN_138; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_140 = 8'h49 == iteration[7:0] ? io_dataIn_73 : _GEN_139; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_141 = 8'h4a == iteration[7:0] ? io_dataIn_74 : _GEN_140; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_142 = 8'h4b == iteration[7:0] ? io_dataIn_75 : _GEN_141; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_143 = 8'h4c == iteration[7:0] ? io_dataIn_76 : _GEN_142; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_144 = 8'h4d == iteration[7:0] ? io_dataIn_77 : _GEN_143; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_145 = 8'h4e == iteration[7:0] ? io_dataIn_78 : _GEN_144; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_146 = 8'h4f == iteration[7:0] ? io_dataIn_79 : _GEN_145; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_147 = 8'h50 == iteration[7:0] ? io_dataIn_80 : _GEN_146; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_148 = 8'h51 == iteration[7:0] ? io_dataIn_81 : _GEN_147; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_149 = 8'h52 == iteration[7:0] ? io_dataIn_82 : _GEN_148; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_150 = 8'h53 == iteration[7:0] ? io_dataIn_83 : _GEN_149; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_151 = 8'h54 == iteration[7:0] ? io_dataIn_84 : _GEN_150; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_152 = 8'h55 == iteration[7:0] ? io_dataIn_85 : _GEN_151; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_153 = 8'h56 == iteration[7:0] ? io_dataIn_86 : _GEN_152; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_154 = 8'h57 == iteration[7:0] ? io_dataIn_87 : _GEN_153; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_155 = 8'h58 == iteration[7:0] ? io_dataIn_88 : _GEN_154; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_156 = 8'h59 == iteration[7:0] ? io_dataIn_89 : _GEN_155; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_157 = 8'h5a == iteration[7:0] ? io_dataIn_90 : _GEN_156; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_158 = 8'h5b == iteration[7:0] ? io_dataIn_91 : _GEN_157; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_159 = 8'h5c == iteration[7:0] ? io_dataIn_92 : _GEN_158; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_160 = 8'h5d == iteration[7:0] ? io_dataIn_93 : _GEN_159; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_161 = 8'h5e == iteration[7:0] ? io_dataIn_94 : _GEN_160; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_162 = 8'h5f == iteration[7:0] ? io_dataIn_95 : _GEN_161; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_163 = 8'h60 == iteration[7:0] ? io_dataIn_96 : _GEN_162; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_164 = 8'h61 == iteration[7:0] ? io_dataIn_97 : _GEN_163; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_165 = 8'h62 == iteration[7:0] ? io_dataIn_98 : _GEN_164; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_166 = 8'h63 == iteration[7:0] ? io_dataIn_99 : _GEN_165; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_167 = 8'h64 == iteration[7:0] ? io_dataIn_100 : _GEN_166; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_168 = 8'h65 == iteration[7:0] ? io_dataIn_101 : _GEN_167; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_169 = 8'h66 == iteration[7:0] ? io_dataIn_102 : _GEN_168; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_170 = 8'h67 == iteration[7:0] ? io_dataIn_103 : _GEN_169; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_171 = 8'h68 == iteration[7:0] ? io_dataIn_104 : _GEN_170; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_172 = 8'h69 == iteration[7:0] ? io_dataIn_105 : _GEN_171; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_173 = 8'h6a == iteration[7:0] ? io_dataIn_106 : _GEN_172; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_174 = 8'h6b == iteration[7:0] ? io_dataIn_107 : _GEN_173; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_175 = 8'h6c == iteration[7:0] ? io_dataIn_108 : _GEN_174; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_176 = 8'h6d == iteration[7:0] ? io_dataIn_109 : _GEN_175; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_177 = 8'h6e == iteration[7:0] ? io_dataIn_110 : _GEN_176; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_178 = 8'h6f == iteration[7:0] ? io_dataIn_111 : _GEN_177; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_179 = 8'h70 == iteration[7:0] ? io_dataIn_112 : _GEN_178; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_180 = 8'h71 == iteration[7:0] ? io_dataIn_113 : _GEN_179; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_181 = 8'h72 == iteration[7:0] ? io_dataIn_114 : _GEN_180; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_182 = 8'h73 == iteration[7:0] ? io_dataIn_115 : _GEN_181; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_183 = 8'h74 == iteration[7:0] ? io_dataIn_116 : _GEN_182; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_184 = 8'h75 == iteration[7:0] ? io_dataIn_117 : _GEN_183; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_185 = 8'h76 == iteration[7:0] ? io_dataIn_118 : _GEN_184; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_186 = 8'h77 == iteration[7:0] ? io_dataIn_119 : _GEN_185; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_187 = 8'h78 == iteration[7:0] ? io_dataIn_120 : _GEN_186; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_188 = 8'h79 == iteration[7:0] ? io_dataIn_121 : _GEN_187; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_189 = 8'h7a == iteration[7:0] ? io_dataIn_122 : _GEN_188; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_190 = 8'h7b == iteration[7:0] ? io_dataIn_123 : _GEN_189; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_191 = 8'h7c == iteration[7:0] ? io_dataIn_124 : _GEN_190; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_192 = 8'h7d == iteration[7:0] ? io_dataIn_125 : _GEN_191; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_193 = 8'h7e == iteration[7:0] ? io_dataIn_126 : _GEN_192; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_194 = 8'h7f == iteration[7:0] ? io_dataIn_127 : _GEN_193; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_195 = 8'h80 == iteration[7:0] ? io_dataIn_128 : _GEN_194; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_196 = 8'h81 == iteration[7:0] ? io_dataIn_129 : _GEN_195; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_197 = 8'h82 == iteration[7:0] ? io_dataIn_130 : _GEN_196; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_198 = 8'h83 == iteration[7:0] ? io_dataIn_131 : _GEN_197; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_199 = 8'h84 == iteration[7:0] ? io_dataIn_132 : _GEN_198; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_200 = 8'h85 == iteration[7:0] ? io_dataIn_133 : _GEN_199; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_201 = 8'h86 == iteration[7:0] ? io_dataIn_134 : _GEN_200; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_202 = 8'h87 == iteration[7:0] ? io_dataIn_135 : _GEN_201; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_203 = 8'h88 == iteration[7:0] ? io_dataIn_136 : _GEN_202; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_204 = 8'h89 == iteration[7:0] ? io_dataIn_137 : _GEN_203; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_205 = 8'h8a == iteration[7:0] ? io_dataIn_138 : _GEN_204; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_206 = 8'h8b == iteration[7:0] ? io_dataIn_139 : _GEN_205; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_207 = 8'h8c == iteration[7:0] ? io_dataIn_140 : _GEN_206; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_208 = 8'h8d == iteration[7:0] ? io_dataIn_141 : _GEN_207; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_209 = 8'h8e == iteration[7:0] ? io_dataIn_142 : _GEN_208; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_210 = 8'h8f == iteration[7:0] ? io_dataIn_143 : _GEN_209; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_211 = 8'h90 == iteration[7:0] ? io_dataIn_144 : _GEN_210; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_212 = 8'h91 == iteration[7:0] ? io_dataIn_145 : _GEN_211; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_213 = 8'h92 == iteration[7:0] ? io_dataIn_146 : _GEN_212; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_214 = 8'h93 == iteration[7:0] ? io_dataIn_147 : _GEN_213; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_215 = 8'h94 == iteration[7:0] ? io_dataIn_148 : _GEN_214; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_216 = 8'h95 == iteration[7:0] ? io_dataIn_149 : _GEN_215; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_217 = 8'h96 == iteration[7:0] ? io_dataIn_150 : _GEN_216; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_218 = 8'h97 == iteration[7:0] ? io_dataIn_151 : _GEN_217; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_219 = 8'h98 == iteration[7:0] ? io_dataIn_152 : _GEN_218; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_220 = 8'h99 == iteration[7:0] ? io_dataIn_153 : _GEN_219; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_221 = 8'h9a == iteration[7:0] ? io_dataIn_154 : _GEN_220; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_222 = 8'h9b == iteration[7:0] ? io_dataIn_155 : _GEN_221; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_223 = 8'h9c == iteration[7:0] ? io_dataIn_156 : _GEN_222; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_224 = 8'h9d == iteration[7:0] ? io_dataIn_157 : _GEN_223; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_225 = 8'h9e == iteration[7:0] ? io_dataIn_158 : _GEN_224; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_226 = 8'h9f == iteration[7:0] ? io_dataIn_159 : _GEN_225; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_227 = 8'ha0 == iteration[7:0] ? io_dataIn_160 : _GEN_226; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_228 = 8'ha1 == iteration[7:0] ? io_dataIn_161 : _GEN_227; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_229 = 8'ha2 == iteration[7:0] ? io_dataIn_162 : _GEN_228; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_230 = 8'ha3 == iteration[7:0] ? io_dataIn_163 : _GEN_229; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_231 = 8'ha4 == iteration[7:0] ? io_dataIn_164 : _GEN_230; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_232 = 8'ha5 == iteration[7:0] ? io_dataIn_165 : _GEN_231; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_233 = 8'ha6 == iteration[7:0] ? io_dataIn_166 : _GEN_232; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_234 = 8'ha7 == iteration[7:0] ? io_dataIn_167 : _GEN_233; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_235 = 8'ha8 == iteration[7:0] ? io_dataIn_168 : _GEN_234; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_236 = 8'ha9 == iteration[7:0] ? io_dataIn_169 : _GEN_235; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_237 = 8'haa == iteration[7:0] ? io_dataIn_170 : _GEN_236; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_238 = 8'hab == iteration[7:0] ? io_dataIn_171 : _GEN_237; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_239 = 8'hac == iteration[7:0] ? io_dataIn_172 : _GEN_238; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_240 = 8'had == iteration[7:0] ? io_dataIn_173 : _GEN_239; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_241 = 8'hae == iteration[7:0] ? io_dataIn_174 : _GEN_240; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_242 = 8'haf == iteration[7:0] ? io_dataIn_175 : _GEN_241; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_243 = 8'hb0 == iteration[7:0] ? io_dataIn_176 : _GEN_242; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_244 = 8'hb1 == iteration[7:0] ? io_dataIn_177 : _GEN_243; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_245 = 8'hb2 == iteration[7:0] ? io_dataIn_178 : _GEN_244; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_246 = 8'hb3 == iteration[7:0] ? io_dataIn_179 : _GEN_245; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_247 = 8'hb4 == iteration[7:0] ? io_dataIn_180 : _GEN_246; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_248 = 8'hb5 == iteration[7:0] ? io_dataIn_181 : _GEN_247; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_249 = 8'hb6 == iteration[7:0] ? io_dataIn_182 : _GEN_248; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_250 = 8'hb7 == iteration[7:0] ? io_dataIn_183 : _GEN_249; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_251 = 8'hb8 == iteration[7:0] ? io_dataIn_184 : _GEN_250; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_252 = 8'hb9 == iteration[7:0] ? io_dataIn_185 : _GEN_251; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_253 = 8'hba == iteration[7:0] ? io_dataIn_186 : _GEN_252; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_254 = 8'hbb == iteration[7:0] ? io_dataIn_187 : _GEN_253; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_255 = 8'hbc == iteration[7:0] ? io_dataIn_188 : _GEN_254; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_256 = 8'hbd == iteration[7:0] ? io_dataIn_189 : _GEN_255; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_257 = 8'hbe == iteration[7:0] ? io_dataIn_190 : _GEN_256; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_258 = 8'hbf == iteration[7:0] ? io_dataIn_191 : _GEN_257; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_259 = 8'hc0 == iteration[7:0] ? io_dataIn_192 : _GEN_258; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_260 = 8'hc1 == iteration[7:0] ? io_dataIn_193 : _GEN_259; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_261 = 8'hc2 == iteration[7:0] ? io_dataIn_194 : _GEN_260; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_262 = 8'hc3 == iteration[7:0] ? io_dataIn_195 : _GEN_261; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_263 = 8'hc4 == iteration[7:0] ? io_dataIn_196 : _GEN_262; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_264 = 8'hc5 == iteration[7:0] ? io_dataIn_197 : _GEN_263; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_265 = 8'hc6 == iteration[7:0] ? io_dataIn_198 : _GEN_264; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_266 = 8'hc7 == iteration[7:0] ? io_dataIn_199 : _GEN_265; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_267 = 8'hc8 == iteration[7:0] ? io_dataIn_200 : _GEN_266; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_268 = 8'hc9 == iteration[7:0] ? io_dataIn_201 : _GEN_267; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_269 = 8'hca == iteration[7:0] ? io_dataIn_202 : _GEN_268; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_270 = 8'hcb == iteration[7:0] ? io_dataIn_203 : _GEN_269; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_271 = 8'hcc == iteration[7:0] ? io_dataIn_204 : _GEN_270; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_272 = 8'hcd == iteration[7:0] ? io_dataIn_205 : _GEN_271; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_273 = 8'hce == iteration[7:0] ? io_dataIn_206 : _GEN_272; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_274 = 8'hcf == iteration[7:0] ? io_dataIn_207 : _GEN_273; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_275 = 8'hd0 == iteration[7:0] ? io_dataIn_208 : _GEN_274; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_276 = 8'hd1 == iteration[7:0] ? io_dataIn_209 : _GEN_275; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_277 = 8'hd2 == iteration[7:0] ? io_dataIn_210 : _GEN_276; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_278 = 8'hd3 == iteration[7:0] ? io_dataIn_211 : _GEN_277; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_279 = 8'hd4 == iteration[7:0] ? io_dataIn_212 : _GEN_278; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_280 = 8'hd5 == iteration[7:0] ? io_dataIn_213 : _GEN_279; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_281 = 8'hd6 == iteration[7:0] ? io_dataIn_214 : _GEN_280; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_282 = 8'hd7 == iteration[7:0] ? io_dataIn_215 : _GEN_281; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_283 = 8'hd8 == iteration[7:0] ? io_dataIn_216 : _GEN_282; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_284 = 8'hd9 == iteration[7:0] ? io_dataIn_217 : _GEN_283; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_285 = 8'hda == iteration[7:0] ? io_dataIn_218 : _GEN_284; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_286 = 8'hdb == iteration[7:0] ? io_dataIn_219 : _GEN_285; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_287 = 8'hdc == iteration[7:0] ? io_dataIn_220 : _GEN_286; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_288 = 8'hdd == iteration[7:0] ? io_dataIn_221 : _GEN_287; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_289 = 8'hde == iteration[7:0] ? io_dataIn_222 : _GEN_288; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_290 = 8'hdf == iteration[7:0] ? io_dataIn_223 : _GEN_289; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_291 = 8'he0 == iteration[7:0] ? io_dataIn_224 : _GEN_290; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_292 = 8'he1 == iteration[7:0] ? io_dataIn_225 : _GEN_291; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_293 = 8'he2 == iteration[7:0] ? io_dataIn_226 : _GEN_292; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_294 = 8'he3 == iteration[7:0] ? io_dataIn_227 : _GEN_293; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_295 = 8'he4 == iteration[7:0] ? io_dataIn_228 : _GEN_294; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_296 = 8'he5 == iteration[7:0] ? io_dataIn_229 : _GEN_295; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_297 = 8'he6 == iteration[7:0] ? io_dataIn_230 : _GEN_296; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_298 = 8'he7 == iteration[7:0] ? io_dataIn_231 : _GEN_297; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_299 = 8'he8 == iteration[7:0] ? io_dataIn_232 : _GEN_298; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_300 = 8'he9 == iteration[7:0] ? io_dataIn_233 : _GEN_299; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_301 = 8'hea == iteration[7:0] ? io_dataIn_234 : _GEN_300; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_302 = 8'heb == iteration[7:0] ? io_dataIn_235 : _GEN_301; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_303 = 8'hec == iteration[7:0] ? io_dataIn_236 : _GEN_302; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_304 = 8'hed == iteration[7:0] ? io_dataIn_237 : _GEN_303; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_305 = 8'hee == iteration[7:0] ? io_dataIn_238 : _GEN_304; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_306 = 8'hef == iteration[7:0] ? io_dataIn_239 : _GEN_305; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_307 = 8'hf0 == iteration[7:0] ? io_dataIn_240 : _GEN_306; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_308 = 8'hf1 == iteration[7:0] ? io_dataIn_241 : _GEN_307; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_309 = 8'hf2 == iteration[7:0] ? io_dataIn_242 : _GEN_308; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_310 = 8'hf3 == iteration[7:0] ? io_dataIn_243 : _GEN_309; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_311 = 8'hf4 == iteration[7:0] ? io_dataIn_244 : _GEN_310; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_312 = 8'hf5 == iteration[7:0] ? io_dataIn_245 : _GEN_311; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_313 = 8'hf6 == iteration[7:0] ? io_dataIn_246 : _GEN_312; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_314 = 8'hf7 == iteration[7:0] ? io_dataIn_247 : _GEN_313; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_315 = 8'hf8 == iteration[7:0] ? io_dataIn_248 : _GEN_314; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_316 = 8'hf9 == iteration[7:0] ? io_dataIn_249 : _GEN_315; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_317 = 8'hfa == iteration[7:0] ? io_dataIn_250 : _GEN_316; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_318 = 8'hfb == iteration[7:0] ? io_dataIn_251 : _GEN_317; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_319 = 8'hfc == iteration[7:0] ? io_dataIn_252 : _GEN_318; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_320 = 8'hfd == iteration[7:0] ? io_dataIn_253 : _GEN_319; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_321 = 8'hfe == iteration[7:0] ? io_dataIn_254 : _GEN_320; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_322 = 8'hff == iteration[7:0] ? io_dataIn_255 : _GEN_321; // @[characterFrequencySort.scala 67:24]
  wire [12:0] _GEN_323 = _T_6 ? _GEN_322 : 13'h0; // @[characterFrequencySort.scala 66:57]
  wire  _T_50 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_51 = iteration == 9'h0; // @[characterFrequencySort.scala 142:22]
  wire [12:0] _GEN_458 = _T_51 ? escapeFrequency : 13'h0; // @[characterFrequencySort.scala 142:31]
  wire [12:0] _GEN_589 = _T_50 ? _GEN_458 : 13'h0; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_721 = _T_4 ? _GEN_323 : _GEN_589; // @[Conditional.scala 39:67]
  wire [12:0] frequencyInput = _T ? 13'h0 : _GEN_721; // @[Conditional.scala 40:58]
  wire  _T_8 = frequencyInput > sortedFrequency_0; // @[characterFrequencySort.scala 75:27]
  wire  _T_9 = sortedFrequencyTemp_0 > sortedFrequency_1; // @[characterFrequencySort.scala 88:49]
  wire  _T_10 = sortedFrequencyTemp_1 > sortedFrequency_2; // @[characterFrequencySort.scala 88:49]
  wire  _T_11 = sortedFrequencyTemp_2 > sortedFrequency_3; // @[characterFrequencySort.scala 88:49]
  wire  _T_12 = sortedFrequencyTemp_3 > sortedFrequency_4; // @[characterFrequencySort.scala 88:49]
  wire  _T_13 = sortedFrequencyTemp_4 > sortedFrequency_5; // @[characterFrequencySort.scala 88:49]
  wire  _T_14 = sortedFrequencyTemp_5 > sortedFrequency_6; // @[characterFrequencySort.scala 88:49]
  wire  _T_15 = sortedFrequencyTemp_6 > sortedFrequency_7; // @[characterFrequencySort.scala 88:49]
  wire  _T_16 = sortedFrequencyTemp_7 > sortedFrequency_8; // @[characterFrequencySort.scala 88:49]
  wire  _T_17 = sortedFrequencyTemp_8 > sortedFrequency_9; // @[characterFrequencySort.scala 88:49]
  wire  _T_18 = sortedFrequencyTemp_9 > sortedFrequency_10; // @[characterFrequencySort.scala 88:49]
  wire  _T_19 = sortedFrequencyTemp_10 > sortedFrequency_11; // @[characterFrequencySort.scala 88:49]
  wire  _T_20 = sortedFrequencyTemp_11 > sortedFrequency_12; // @[characterFrequencySort.scala 88:49]
  wire  _T_21 = sortedFrequencyTemp_12 > sortedFrequency_13; // @[characterFrequencySort.scala 88:49]
  wire  _T_22 = sortedFrequencyTemp_13 > sortedFrequency_14; // @[characterFrequencySort.scala 88:49]
  wire  _T_23 = sortedFrequencyTemp_14 > sortedFrequency_15; // @[characterFrequencySort.scala 88:49]
  wire  _T_24 = sortedFrequencyTemp_15 > sortedFrequency_16; // @[characterFrequencySort.scala 88:49]
  wire  _T_25 = sortedFrequencyTemp_16 > sortedFrequency_17; // @[characterFrequencySort.scala 88:49]
  wire  _T_26 = sortedFrequencyTemp_17 > sortedFrequency_18; // @[characterFrequencySort.scala 88:49]
  wire  _T_27 = sortedFrequencyTemp_18 > sortedFrequency_19; // @[characterFrequencySort.scala 88:49]
  wire  _T_28 = sortedFrequencyTemp_19 > sortedFrequency_20; // @[characterFrequencySort.scala 88:49]
  wire  _T_29 = sortedFrequencyTemp_20 > sortedFrequency_21; // @[characterFrequencySort.scala 88:49]
  wire  _T_30 = sortedFrequencyTemp_21 > sortedFrequency_22; // @[characterFrequencySort.scala 88:49]
  wire  _T_31 = sortedFrequencyTemp_22 > sortedFrequency_23; // @[characterFrequencySort.scala 88:49]
  wire  _T_32 = sortedFrequencyTemp_23 > sortedFrequency_24; // @[characterFrequencySort.scala 88:49]
  wire  _T_33 = sortedFrequencyTemp_24 > sortedFrequency_25; // @[characterFrequencySort.scala 88:49]
  wire  _T_34 = sortedFrequencyTemp_25 > sortedFrequency_26; // @[characterFrequencySort.scala 88:49]
  wire  _T_35 = sortedFrequencyTemp_26 > sortedFrequency_27; // @[characterFrequencySort.scala 88:49]
  wire  _T_36 = sortedFrequencyTemp_27 > sortedFrequency_28; // @[characterFrequencySort.scala 88:49]
  wire  _T_37 = sortedFrequencyTemp_28 > sortedFrequency_29; // @[characterFrequencySort.scala 88:49]
  wire  _T_38 = sortedFrequencyTemp_29 > sortedFrequency_30; // @[characterFrequencySort.scala 88:49]
  wire  _T_39 = sortedFrequencyTemp_30 > sortedFrequency_31; // @[characterFrequencySort.scala 101:67]
  wire [12:0] _T_41 = escapeFrequency + sortedFrequency_31; // @[characterFrequencySort.scala 105:44]
  wire [12:0] _T_43 = escapeFrequency + sortedFrequencyTemp_30; // @[characterFrequencySort.scala 115:44]
  wire [8:0] _T_45 = iteration + 9'h1; // @[characterFrequencySort.scala 120:30]
  wire  _T_46 = iteration == 9'h11f; // @[characterFrequencySort.scala 121:22]
  wire  _T_47 = escapeFrequency > 13'h0; // @[characterFrequencySort.scala 124:30]
  wire  _T_86 = iteration == 9'h1f; // @[characterFrequencySort.scala 177:22]
  assign io_sortedFrequency_0 = sortedFrequency_0; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_1 = sortedFrequency_1; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_2 = sortedFrequency_2; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_3 = sortedFrequency_3; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_4 = sortedFrequency_4; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_5 = sortedFrequency_5; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_6 = sortedFrequency_6; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_7 = sortedFrequency_7; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_8 = sortedFrequency_8; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_9 = sortedFrequency_9; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_10 = sortedFrequency_10; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_11 = sortedFrequency_11; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_12 = sortedFrequency_12; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_13 = sortedFrequency_13; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_14 = sortedFrequency_14; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_15 = sortedFrequency_15; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_16 = sortedFrequency_16; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_17 = sortedFrequency_17; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_18 = sortedFrequency_18; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_19 = sortedFrequency_19; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_20 = sortedFrequency_20; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_21 = sortedFrequency_21; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_22 = sortedFrequency_22; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_23 = sortedFrequency_23; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_24 = sortedFrequency_24; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_25 = sortedFrequency_25; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_26 = sortedFrequency_26; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_27 = sortedFrequency_27; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_28 = sortedFrequency_28; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_29 = sortedFrequency_29; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_30 = sortedFrequency_30; // @[characterFrequencySort.scala 184:22]
  assign io_sortedFrequency_31 = sortedFrequency_31; // @[characterFrequencySort.scala 184:22]
  assign io_sortedCharacter_0 = sortedCharacter_0; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_1 = sortedCharacter_1; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_2 = sortedCharacter_2; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_3 = sortedCharacter_3; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_4 = sortedCharacter_4; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_5 = sortedCharacter_5; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_6 = sortedCharacter_6; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_7 = sortedCharacter_7; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_8 = sortedCharacter_8; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_9 = sortedCharacter_9; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_10 = sortedCharacter_10; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_11 = sortedCharacter_11; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_12 = sortedCharacter_12; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_13 = sortedCharacter_13; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_14 = sortedCharacter_14; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_15 = sortedCharacter_15; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_16 = sortedCharacter_16; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_17 = sortedCharacter_17; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_18 = sortedCharacter_18; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_19 = sortedCharacter_19; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_20 = sortedCharacter_20; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_21 = sortedCharacter_21; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_22 = sortedCharacter_22; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_23 = sortedCharacter_23; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_24 = sortedCharacter_24; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_25 = sortedCharacter_25; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_26 = sortedCharacter_26; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_27 = sortedCharacter_27; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_28 = sortedCharacter_28; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_29 = sortedCharacter_29; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_30 = sortedCharacter_30; // @[characterFrequencySort.scala 185:22]
  assign io_sortedCharacter_31 = sortedCharacter_31; // @[characterFrequencySort.scala 185:22]
  assign io_finished = state == 2'h0; // @[characterFrequencySort.scala 183:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  iteration = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  sortedFrequency_0 = _RAND_2[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  sortedFrequency_1 = _RAND_3[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  sortedFrequency_2 = _RAND_4[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sortedFrequency_3 = _RAND_5[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sortedFrequency_4 = _RAND_6[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sortedFrequency_5 = _RAND_7[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sortedFrequency_6 = _RAND_8[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  sortedFrequency_7 = _RAND_9[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  sortedFrequency_8 = _RAND_10[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  sortedFrequency_9 = _RAND_11[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  sortedFrequency_10 = _RAND_12[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  sortedFrequency_11 = _RAND_13[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  sortedFrequency_12 = _RAND_14[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  sortedFrequency_13 = _RAND_15[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  sortedFrequency_14 = _RAND_16[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  sortedFrequency_15 = _RAND_17[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  sortedFrequency_16 = _RAND_18[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  sortedFrequency_17 = _RAND_19[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  sortedFrequency_18 = _RAND_20[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  sortedFrequency_19 = _RAND_21[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  sortedFrequency_20 = _RAND_22[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  sortedFrequency_21 = _RAND_23[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  sortedFrequency_22 = _RAND_24[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  sortedFrequency_23 = _RAND_25[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  sortedFrequency_24 = _RAND_26[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  sortedFrequency_25 = _RAND_27[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  sortedFrequency_26 = _RAND_28[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  sortedFrequency_27 = _RAND_29[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  sortedFrequency_28 = _RAND_30[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  sortedFrequency_29 = _RAND_31[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  sortedFrequency_30 = _RAND_32[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  sortedFrequency_31 = _RAND_33[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  sortedCharacter_0 = _RAND_34[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  sortedCharacter_1 = _RAND_35[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  sortedCharacter_2 = _RAND_36[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  sortedCharacter_3 = _RAND_37[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  sortedCharacter_4 = _RAND_38[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  sortedCharacter_5 = _RAND_39[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  sortedCharacter_6 = _RAND_40[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  sortedCharacter_7 = _RAND_41[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  sortedCharacter_8 = _RAND_42[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  sortedCharacter_9 = _RAND_43[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  sortedCharacter_10 = _RAND_44[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  sortedCharacter_11 = _RAND_45[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  sortedCharacter_12 = _RAND_46[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  sortedCharacter_13 = _RAND_47[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  sortedCharacter_14 = _RAND_48[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  sortedCharacter_15 = _RAND_49[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  sortedCharacter_16 = _RAND_50[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  sortedCharacter_17 = _RAND_51[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  sortedCharacter_18 = _RAND_52[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  sortedCharacter_19 = _RAND_53[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  sortedCharacter_20 = _RAND_54[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  sortedCharacter_21 = _RAND_55[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  sortedCharacter_22 = _RAND_56[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  sortedCharacter_23 = _RAND_57[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  sortedCharacter_24 = _RAND_58[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  sortedCharacter_25 = _RAND_59[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  sortedCharacter_26 = _RAND_60[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  sortedCharacter_27 = _RAND_61[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  sortedCharacter_28 = _RAND_62[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  sortedCharacter_29 = _RAND_63[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  sortedCharacter_30 = _RAND_64[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  sortedCharacter_31 = _RAND_65[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  sortedFrequencyTemp_0 = _RAND_66[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  sortedFrequencyTemp_1 = _RAND_67[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  sortedFrequencyTemp_2 = _RAND_68[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  sortedFrequencyTemp_3 = _RAND_69[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  sortedFrequencyTemp_4 = _RAND_70[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  sortedFrequencyTemp_5 = _RAND_71[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  sortedFrequencyTemp_6 = _RAND_72[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  sortedFrequencyTemp_7 = _RAND_73[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  sortedFrequencyTemp_8 = _RAND_74[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  sortedFrequencyTemp_9 = _RAND_75[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  sortedFrequencyTemp_10 = _RAND_76[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  sortedFrequencyTemp_11 = _RAND_77[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  sortedFrequencyTemp_12 = _RAND_78[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  sortedFrequencyTemp_13 = _RAND_79[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  sortedFrequencyTemp_14 = _RAND_80[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  sortedFrequencyTemp_15 = _RAND_81[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  sortedFrequencyTemp_16 = _RAND_82[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  sortedFrequencyTemp_17 = _RAND_83[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  sortedFrequencyTemp_18 = _RAND_84[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  sortedFrequencyTemp_19 = _RAND_85[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  sortedFrequencyTemp_20 = _RAND_86[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  sortedFrequencyTemp_21 = _RAND_87[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  sortedFrequencyTemp_22 = _RAND_88[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  sortedFrequencyTemp_23 = _RAND_89[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  sortedFrequencyTemp_24 = _RAND_90[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  sortedFrequencyTemp_25 = _RAND_91[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  sortedFrequencyTemp_26 = _RAND_92[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  sortedFrequencyTemp_27 = _RAND_93[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  sortedFrequencyTemp_28 = _RAND_94[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  sortedFrequencyTemp_29 = _RAND_95[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  sortedFrequencyTemp_30 = _RAND_96[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  sortedCharacterTemp_0 = _RAND_97[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  sortedCharacterTemp_1 = _RAND_98[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  sortedCharacterTemp_2 = _RAND_99[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  sortedCharacterTemp_3 = _RAND_100[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  sortedCharacterTemp_4 = _RAND_101[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  sortedCharacterTemp_5 = _RAND_102[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  sortedCharacterTemp_6 = _RAND_103[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  sortedCharacterTemp_7 = _RAND_104[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  sortedCharacterTemp_8 = _RAND_105[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  sortedCharacterTemp_9 = _RAND_106[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  sortedCharacterTemp_10 = _RAND_107[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  sortedCharacterTemp_11 = _RAND_108[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  sortedCharacterTemp_12 = _RAND_109[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  sortedCharacterTemp_13 = _RAND_110[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  sortedCharacterTemp_14 = _RAND_111[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  sortedCharacterTemp_15 = _RAND_112[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  sortedCharacterTemp_16 = _RAND_113[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  sortedCharacterTemp_17 = _RAND_114[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  sortedCharacterTemp_18 = _RAND_115[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  sortedCharacterTemp_19 = _RAND_116[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  sortedCharacterTemp_20 = _RAND_117[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  sortedCharacterTemp_21 = _RAND_118[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  sortedCharacterTemp_22 = _RAND_119[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  sortedCharacterTemp_23 = _RAND_120[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  sortedCharacterTemp_24 = _RAND_121[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  sortedCharacterTemp_25 = _RAND_122[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  sortedCharacterTemp_26 = _RAND_123[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  sortedCharacterTemp_27 = _RAND_124[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  sortedCharacterTemp_28 = _RAND_125[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  sortedCharacterTemp_29 = _RAND_126[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  sortedCharacterTemp_30 = _RAND_127[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  escapeFrequency = _RAND_128[12:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T) begin
      if (io_start) begin
        state <= 2'h1;
      end
    end else if (_T_4) begin
      if (_T_46) begin
        if (_T_47) begin
          state <= 2'h2;
        end else begin
          state <= 2'h0;
        end
      end
    end else if (_T_50) begin
      if (_T_86) begin
        state <= 2'h0;
      end
    end
    if (_T) begin
      if (io_start) begin
        iteration <= 9'h0;
      end
    end else if (_T_4) begin
      if (_T_46) begin
        if (_T_47) begin
          iteration <= 9'h0;
        end else begin
          iteration <= _T_45;
        end
      end else begin
        iteration <= _T_45;
      end
    end else if (_T_50) begin
      iteration <= _T_45;
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_0 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_8) begin
        if (_T) begin
          sortedFrequency_0 <= 13'h0;
        end else if (_T_4) begin
          if (_T_6) begin
            if (8'hff == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_255;
            end else if (8'hfe == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_254;
            end else if (8'hfd == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_253;
            end else if (8'hfc == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_252;
            end else if (8'hfb == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_251;
            end else if (8'hfa == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_250;
            end else if (8'hf9 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_249;
            end else if (8'hf8 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_248;
            end else if (8'hf7 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_247;
            end else if (8'hf6 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_246;
            end else if (8'hf5 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_245;
            end else if (8'hf4 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_244;
            end else if (8'hf3 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_243;
            end else if (8'hf2 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_242;
            end else if (8'hf1 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_241;
            end else if (8'hf0 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_240;
            end else if (8'hef == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_239;
            end else if (8'hee == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_238;
            end else if (8'hed == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_237;
            end else if (8'hec == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_236;
            end else if (8'heb == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_235;
            end else if (8'hea == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_234;
            end else if (8'he9 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_233;
            end else if (8'he8 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_232;
            end else if (8'he7 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_231;
            end else if (8'he6 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_230;
            end else if (8'he5 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_229;
            end else if (8'he4 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_228;
            end else if (8'he3 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_227;
            end else if (8'he2 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_226;
            end else if (8'he1 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_225;
            end else if (8'he0 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_224;
            end else if (8'hdf == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_223;
            end else if (8'hde == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_222;
            end else if (8'hdd == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_221;
            end else if (8'hdc == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_220;
            end else if (8'hdb == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_219;
            end else if (8'hda == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_218;
            end else if (8'hd9 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_217;
            end else if (8'hd8 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_216;
            end else if (8'hd7 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_215;
            end else if (8'hd6 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_214;
            end else if (8'hd5 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_213;
            end else if (8'hd4 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_212;
            end else if (8'hd3 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_211;
            end else if (8'hd2 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_210;
            end else if (8'hd1 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_209;
            end else if (8'hd0 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_208;
            end else if (8'hcf == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_207;
            end else if (8'hce == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_206;
            end else if (8'hcd == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_205;
            end else if (8'hcc == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_204;
            end else if (8'hcb == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_203;
            end else if (8'hca == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_202;
            end else if (8'hc9 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_201;
            end else if (8'hc8 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_200;
            end else if (8'hc7 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_199;
            end else if (8'hc6 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_198;
            end else if (8'hc5 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_197;
            end else if (8'hc4 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_196;
            end else if (8'hc3 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_195;
            end else if (8'hc2 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_194;
            end else if (8'hc1 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_193;
            end else if (8'hc0 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_192;
            end else if (8'hbf == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_191;
            end else if (8'hbe == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_190;
            end else if (8'hbd == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_189;
            end else if (8'hbc == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_188;
            end else if (8'hbb == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_187;
            end else if (8'hba == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_186;
            end else if (8'hb9 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_185;
            end else if (8'hb8 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_184;
            end else if (8'hb7 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_183;
            end else if (8'hb6 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_182;
            end else if (8'hb5 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_181;
            end else if (8'hb4 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_180;
            end else if (8'hb3 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_179;
            end else if (8'hb2 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_178;
            end else if (8'hb1 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_177;
            end else if (8'hb0 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_176;
            end else if (8'haf == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_175;
            end else if (8'hae == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_174;
            end else if (8'had == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_173;
            end else if (8'hac == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_172;
            end else if (8'hab == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_171;
            end else if (8'haa == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_170;
            end else if (8'ha9 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_169;
            end else if (8'ha8 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_168;
            end else if (8'ha7 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_167;
            end else if (8'ha6 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_166;
            end else if (8'ha5 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_165;
            end else if (8'ha4 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_164;
            end else if (8'ha3 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_163;
            end else if (8'ha2 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_162;
            end else if (8'ha1 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_161;
            end else if (8'ha0 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_160;
            end else if (8'h9f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_159;
            end else if (8'h9e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_158;
            end else if (8'h9d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_157;
            end else if (8'h9c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_156;
            end else if (8'h9b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_155;
            end else if (8'h9a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_154;
            end else if (8'h99 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_153;
            end else if (8'h98 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_152;
            end else if (8'h97 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_151;
            end else if (8'h96 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_150;
            end else if (8'h95 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_149;
            end else if (8'h94 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_148;
            end else if (8'h93 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_147;
            end else if (8'h92 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_146;
            end else if (8'h91 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_145;
            end else if (8'h90 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_144;
            end else if (8'h8f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_143;
            end else if (8'h8e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_142;
            end else if (8'h8d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_141;
            end else if (8'h8c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_140;
            end else if (8'h8b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_139;
            end else if (8'h8a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_138;
            end else if (8'h89 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_137;
            end else if (8'h88 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_136;
            end else if (8'h87 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_135;
            end else if (8'h86 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_134;
            end else if (8'h85 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_133;
            end else if (8'h84 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_132;
            end else if (8'h83 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_131;
            end else if (8'h82 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_130;
            end else if (8'h81 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_129;
            end else if (8'h80 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_128;
            end else if (8'h7f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_127;
            end else if (8'h7e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_126;
            end else if (8'h7d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_125;
            end else if (8'h7c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_124;
            end else if (8'h7b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_123;
            end else if (8'h7a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_122;
            end else if (8'h79 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_121;
            end else if (8'h78 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_120;
            end else if (8'h77 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_119;
            end else if (8'h76 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_118;
            end else if (8'h75 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_117;
            end else if (8'h74 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_116;
            end else if (8'h73 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_115;
            end else if (8'h72 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_114;
            end else if (8'h71 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_113;
            end else if (8'h70 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_112;
            end else if (8'h6f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_111;
            end else if (8'h6e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_110;
            end else if (8'h6d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_109;
            end else if (8'h6c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_108;
            end else if (8'h6b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_107;
            end else if (8'h6a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_106;
            end else if (8'h69 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_105;
            end else if (8'h68 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_104;
            end else if (8'h67 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_103;
            end else if (8'h66 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_102;
            end else if (8'h65 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_101;
            end else if (8'h64 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_100;
            end else if (8'h63 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_99;
            end else if (8'h62 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_98;
            end else if (8'h61 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_97;
            end else if (8'h60 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_96;
            end else if (8'h5f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_95;
            end else if (8'h5e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_94;
            end else if (8'h5d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_93;
            end else if (8'h5c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_92;
            end else if (8'h5b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_91;
            end else if (8'h5a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_90;
            end else if (8'h59 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_89;
            end else if (8'h58 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_88;
            end else if (8'h57 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_87;
            end else if (8'h56 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_86;
            end else if (8'h55 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_85;
            end else if (8'h54 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_84;
            end else if (8'h53 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_83;
            end else if (8'h52 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_82;
            end else if (8'h51 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_81;
            end else if (8'h50 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_80;
            end else if (8'h4f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_79;
            end else if (8'h4e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_78;
            end else if (8'h4d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_77;
            end else if (8'h4c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_76;
            end else if (8'h4b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_75;
            end else if (8'h4a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_74;
            end else if (8'h49 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_73;
            end else if (8'h48 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_72;
            end else if (8'h47 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_71;
            end else if (8'h46 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_70;
            end else if (8'h45 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_69;
            end else if (8'h44 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_68;
            end else if (8'h43 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_67;
            end else if (8'h42 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_66;
            end else if (8'h41 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_65;
            end else if (8'h40 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_64;
            end else if (8'h3f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_63;
            end else if (8'h3e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_62;
            end else if (8'h3d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_61;
            end else if (8'h3c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_60;
            end else if (8'h3b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_59;
            end else if (8'h3a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_58;
            end else if (8'h39 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_57;
            end else if (8'h38 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_56;
            end else if (8'h37 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_55;
            end else if (8'h36 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_54;
            end else if (8'h35 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_53;
            end else if (8'h34 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_52;
            end else if (8'h33 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_51;
            end else if (8'h32 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_50;
            end else if (8'h31 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_49;
            end else if (8'h30 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_48;
            end else if (8'h2f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_47;
            end else if (8'h2e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_46;
            end else if (8'h2d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_45;
            end else if (8'h2c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_44;
            end else if (8'h2b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_43;
            end else if (8'h2a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_42;
            end else if (8'h29 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_41;
            end else if (8'h28 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_40;
            end else if (8'h27 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_39;
            end else if (8'h26 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_38;
            end else if (8'h25 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_37;
            end else if (8'h24 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_36;
            end else if (8'h23 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_35;
            end else if (8'h22 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_34;
            end else if (8'h21 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_33;
            end else if (8'h20 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_32;
            end else if (8'h1f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_31;
            end else if (8'h1e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_30;
            end else if (8'h1d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_29;
            end else if (8'h1c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_28;
            end else if (8'h1b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_27;
            end else if (8'h1a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_26;
            end else if (8'h19 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_25;
            end else if (8'h18 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_24;
            end else if (8'h17 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_23;
            end else if (8'h16 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_22;
            end else if (8'h15 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_21;
            end else if (8'h14 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_20;
            end else if (8'h13 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_19;
            end else if (8'h12 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_18;
            end else if (8'h11 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_17;
            end else if (8'h10 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_16;
            end else if (8'hf == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_15;
            end else if (8'he == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_14;
            end else if (8'hd == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_13;
            end else if (8'hc == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_12;
            end else if (8'hb == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_11;
            end else if (8'ha == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_10;
            end else if (8'h9 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_9;
            end else if (8'h8 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_8;
            end else if (8'h7 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_7;
            end else if (8'h6 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_6;
            end else if (8'h5 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_5;
            end else if (8'h4 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_4;
            end else if (8'h3 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_3;
            end else if (8'h2 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_2;
            end else if (8'h1 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_1;
            end else begin
              sortedFrequency_0 <= io_dataIn_0;
            end
          end else begin
            sortedFrequency_0 <= 13'h0;
          end
        end else if (_T_50) begin
          if (_T_51) begin
            sortedFrequency_0 <= escapeFrequency;
          end else begin
            sortedFrequency_0 <= 13'h0;
          end
        end else begin
          sortedFrequency_0 <= 13'h0;
        end
      end
    end else if (_T_50) begin
      if (_T_8) begin
        if (_T) begin
          sortedFrequency_0 <= 13'h0;
        end else if (_T_4) begin
          if (_T_6) begin
            if (8'hff == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_255;
            end else if (8'hfe == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_254;
            end else if (8'hfd == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_253;
            end else if (8'hfc == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_252;
            end else if (8'hfb == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_251;
            end else if (8'hfa == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_250;
            end else if (8'hf9 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_249;
            end else if (8'hf8 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_248;
            end else if (8'hf7 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_247;
            end else if (8'hf6 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_246;
            end else if (8'hf5 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_245;
            end else if (8'hf4 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_244;
            end else if (8'hf3 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_243;
            end else if (8'hf2 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_242;
            end else if (8'hf1 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_241;
            end else if (8'hf0 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_240;
            end else if (8'hef == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_239;
            end else if (8'hee == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_238;
            end else if (8'hed == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_237;
            end else if (8'hec == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_236;
            end else if (8'heb == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_235;
            end else if (8'hea == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_234;
            end else if (8'he9 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_233;
            end else if (8'he8 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_232;
            end else if (8'he7 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_231;
            end else if (8'he6 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_230;
            end else if (8'he5 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_229;
            end else if (8'he4 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_228;
            end else if (8'he3 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_227;
            end else if (8'he2 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_226;
            end else if (8'he1 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_225;
            end else if (8'he0 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_224;
            end else if (8'hdf == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_223;
            end else if (8'hde == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_222;
            end else if (8'hdd == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_221;
            end else if (8'hdc == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_220;
            end else if (8'hdb == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_219;
            end else if (8'hda == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_218;
            end else if (8'hd9 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_217;
            end else if (8'hd8 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_216;
            end else if (8'hd7 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_215;
            end else if (8'hd6 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_214;
            end else if (8'hd5 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_213;
            end else if (8'hd4 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_212;
            end else if (8'hd3 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_211;
            end else if (8'hd2 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_210;
            end else if (8'hd1 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_209;
            end else if (8'hd0 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_208;
            end else if (8'hcf == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_207;
            end else if (8'hce == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_206;
            end else if (8'hcd == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_205;
            end else if (8'hcc == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_204;
            end else if (8'hcb == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_203;
            end else if (8'hca == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_202;
            end else if (8'hc9 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_201;
            end else if (8'hc8 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_200;
            end else if (8'hc7 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_199;
            end else if (8'hc6 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_198;
            end else if (8'hc5 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_197;
            end else if (8'hc4 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_196;
            end else if (8'hc3 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_195;
            end else if (8'hc2 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_194;
            end else if (8'hc1 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_193;
            end else if (8'hc0 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_192;
            end else if (8'hbf == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_191;
            end else if (8'hbe == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_190;
            end else if (8'hbd == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_189;
            end else if (8'hbc == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_188;
            end else if (8'hbb == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_187;
            end else if (8'hba == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_186;
            end else if (8'hb9 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_185;
            end else if (8'hb8 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_184;
            end else if (8'hb7 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_183;
            end else if (8'hb6 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_182;
            end else if (8'hb5 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_181;
            end else if (8'hb4 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_180;
            end else if (8'hb3 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_179;
            end else if (8'hb2 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_178;
            end else if (8'hb1 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_177;
            end else if (8'hb0 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_176;
            end else if (8'haf == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_175;
            end else if (8'hae == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_174;
            end else if (8'had == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_173;
            end else if (8'hac == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_172;
            end else if (8'hab == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_171;
            end else if (8'haa == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_170;
            end else if (8'ha9 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_169;
            end else if (8'ha8 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_168;
            end else if (8'ha7 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_167;
            end else if (8'ha6 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_166;
            end else if (8'ha5 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_165;
            end else if (8'ha4 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_164;
            end else if (8'ha3 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_163;
            end else if (8'ha2 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_162;
            end else if (8'ha1 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_161;
            end else if (8'ha0 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_160;
            end else if (8'h9f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_159;
            end else if (8'h9e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_158;
            end else if (8'h9d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_157;
            end else if (8'h9c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_156;
            end else if (8'h9b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_155;
            end else if (8'h9a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_154;
            end else if (8'h99 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_153;
            end else if (8'h98 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_152;
            end else if (8'h97 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_151;
            end else if (8'h96 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_150;
            end else if (8'h95 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_149;
            end else if (8'h94 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_148;
            end else if (8'h93 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_147;
            end else if (8'h92 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_146;
            end else if (8'h91 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_145;
            end else if (8'h90 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_144;
            end else if (8'h8f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_143;
            end else if (8'h8e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_142;
            end else if (8'h8d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_141;
            end else if (8'h8c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_140;
            end else if (8'h8b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_139;
            end else if (8'h8a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_138;
            end else if (8'h89 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_137;
            end else if (8'h88 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_136;
            end else if (8'h87 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_135;
            end else if (8'h86 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_134;
            end else if (8'h85 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_133;
            end else if (8'h84 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_132;
            end else if (8'h83 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_131;
            end else if (8'h82 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_130;
            end else if (8'h81 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_129;
            end else if (8'h80 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_128;
            end else if (8'h7f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_127;
            end else if (8'h7e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_126;
            end else if (8'h7d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_125;
            end else if (8'h7c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_124;
            end else if (8'h7b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_123;
            end else if (8'h7a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_122;
            end else if (8'h79 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_121;
            end else if (8'h78 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_120;
            end else if (8'h77 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_119;
            end else if (8'h76 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_118;
            end else if (8'h75 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_117;
            end else if (8'h74 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_116;
            end else if (8'h73 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_115;
            end else if (8'h72 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_114;
            end else if (8'h71 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_113;
            end else if (8'h70 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_112;
            end else if (8'h6f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_111;
            end else if (8'h6e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_110;
            end else if (8'h6d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_109;
            end else if (8'h6c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_108;
            end else if (8'h6b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_107;
            end else if (8'h6a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_106;
            end else if (8'h69 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_105;
            end else if (8'h68 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_104;
            end else if (8'h67 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_103;
            end else if (8'h66 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_102;
            end else if (8'h65 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_101;
            end else if (8'h64 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_100;
            end else if (8'h63 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_99;
            end else if (8'h62 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_98;
            end else if (8'h61 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_97;
            end else if (8'h60 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_96;
            end else if (8'h5f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_95;
            end else if (8'h5e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_94;
            end else if (8'h5d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_93;
            end else if (8'h5c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_92;
            end else if (8'h5b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_91;
            end else if (8'h5a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_90;
            end else if (8'h59 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_89;
            end else if (8'h58 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_88;
            end else if (8'h57 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_87;
            end else if (8'h56 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_86;
            end else if (8'h55 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_85;
            end else if (8'h54 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_84;
            end else if (8'h53 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_83;
            end else if (8'h52 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_82;
            end else if (8'h51 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_81;
            end else if (8'h50 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_80;
            end else if (8'h4f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_79;
            end else if (8'h4e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_78;
            end else if (8'h4d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_77;
            end else if (8'h4c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_76;
            end else if (8'h4b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_75;
            end else if (8'h4a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_74;
            end else if (8'h49 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_73;
            end else if (8'h48 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_72;
            end else if (8'h47 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_71;
            end else if (8'h46 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_70;
            end else if (8'h45 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_69;
            end else if (8'h44 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_68;
            end else if (8'h43 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_67;
            end else if (8'h42 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_66;
            end else if (8'h41 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_65;
            end else if (8'h40 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_64;
            end else if (8'h3f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_63;
            end else if (8'h3e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_62;
            end else if (8'h3d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_61;
            end else if (8'h3c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_60;
            end else if (8'h3b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_59;
            end else if (8'h3a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_58;
            end else if (8'h39 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_57;
            end else if (8'h38 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_56;
            end else if (8'h37 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_55;
            end else if (8'h36 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_54;
            end else if (8'h35 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_53;
            end else if (8'h34 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_52;
            end else if (8'h33 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_51;
            end else if (8'h32 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_50;
            end else if (8'h31 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_49;
            end else if (8'h30 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_48;
            end else if (8'h2f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_47;
            end else if (8'h2e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_46;
            end else if (8'h2d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_45;
            end else if (8'h2c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_44;
            end else if (8'h2b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_43;
            end else if (8'h2a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_42;
            end else if (8'h29 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_41;
            end else if (8'h28 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_40;
            end else if (8'h27 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_39;
            end else if (8'h26 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_38;
            end else if (8'h25 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_37;
            end else if (8'h24 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_36;
            end else if (8'h23 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_35;
            end else if (8'h22 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_34;
            end else if (8'h21 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_33;
            end else if (8'h20 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_32;
            end else if (8'h1f == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_31;
            end else if (8'h1e == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_30;
            end else if (8'h1d == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_29;
            end else if (8'h1c == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_28;
            end else if (8'h1b == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_27;
            end else if (8'h1a == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_26;
            end else if (8'h19 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_25;
            end else if (8'h18 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_24;
            end else if (8'h17 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_23;
            end else if (8'h16 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_22;
            end else if (8'h15 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_21;
            end else if (8'h14 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_20;
            end else if (8'h13 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_19;
            end else if (8'h12 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_18;
            end else if (8'h11 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_17;
            end else if (8'h10 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_16;
            end else if (8'hf == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_15;
            end else if (8'he == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_14;
            end else if (8'hd == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_13;
            end else if (8'hc == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_12;
            end else if (8'hb == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_11;
            end else if (8'ha == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_10;
            end else if (8'h9 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_9;
            end else if (8'h8 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_8;
            end else if (8'h7 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_7;
            end else if (8'h6 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_6;
            end else if (8'h5 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_5;
            end else if (8'h4 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_4;
            end else if (8'h3 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_3;
            end else if (8'h2 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_2;
            end else if (8'h1 == iteration[7:0]) begin
              sortedFrequency_0 <= io_dataIn_1;
            end else begin
              sortedFrequency_0 <= io_dataIn_0;
            end
          end else begin
            sortedFrequency_0 <= 13'h0;
          end
        end else if (_T_50) begin
          if (_T_51) begin
            sortedFrequency_0 <= escapeFrequency;
          end else begin
            sortedFrequency_0 <= 13'h0;
          end
        end else begin
          sortedFrequency_0 <= 13'h0;
        end
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_1 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_9) begin
        sortedFrequency_1 <= sortedFrequencyTemp_0;
      end
    end else if (_T_50) begin
      if (_T_9) begin
        sortedFrequency_1 <= sortedFrequencyTemp_0;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_2 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_10) begin
        sortedFrequency_2 <= sortedFrequencyTemp_1;
      end
    end else if (_T_50) begin
      if (_T_10) begin
        sortedFrequency_2 <= sortedFrequencyTemp_1;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_3 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_11) begin
        sortedFrequency_3 <= sortedFrequencyTemp_2;
      end
    end else if (_T_50) begin
      if (_T_11) begin
        sortedFrequency_3 <= sortedFrequencyTemp_2;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_4 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_12) begin
        sortedFrequency_4 <= sortedFrequencyTemp_3;
      end
    end else if (_T_50) begin
      if (_T_12) begin
        sortedFrequency_4 <= sortedFrequencyTemp_3;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_5 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_13) begin
        sortedFrequency_5 <= sortedFrequencyTemp_4;
      end
    end else if (_T_50) begin
      if (_T_13) begin
        sortedFrequency_5 <= sortedFrequencyTemp_4;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_6 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_14) begin
        sortedFrequency_6 <= sortedFrequencyTemp_5;
      end
    end else if (_T_50) begin
      if (_T_14) begin
        sortedFrequency_6 <= sortedFrequencyTemp_5;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_7 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_15) begin
        sortedFrequency_7 <= sortedFrequencyTemp_6;
      end
    end else if (_T_50) begin
      if (_T_15) begin
        sortedFrequency_7 <= sortedFrequencyTemp_6;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_8 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_16) begin
        sortedFrequency_8 <= sortedFrequencyTemp_7;
      end
    end else if (_T_50) begin
      if (_T_16) begin
        sortedFrequency_8 <= sortedFrequencyTemp_7;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_9 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_17) begin
        sortedFrequency_9 <= sortedFrequencyTemp_8;
      end
    end else if (_T_50) begin
      if (_T_17) begin
        sortedFrequency_9 <= sortedFrequencyTemp_8;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_10 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_18) begin
        sortedFrequency_10 <= sortedFrequencyTemp_9;
      end
    end else if (_T_50) begin
      if (_T_18) begin
        sortedFrequency_10 <= sortedFrequencyTemp_9;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_11 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_19) begin
        sortedFrequency_11 <= sortedFrequencyTemp_10;
      end
    end else if (_T_50) begin
      if (_T_19) begin
        sortedFrequency_11 <= sortedFrequencyTemp_10;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_12 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_20) begin
        sortedFrequency_12 <= sortedFrequencyTemp_11;
      end
    end else if (_T_50) begin
      if (_T_20) begin
        sortedFrequency_12 <= sortedFrequencyTemp_11;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_13 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_21) begin
        sortedFrequency_13 <= sortedFrequencyTemp_12;
      end
    end else if (_T_50) begin
      if (_T_21) begin
        sortedFrequency_13 <= sortedFrequencyTemp_12;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_14 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_22) begin
        sortedFrequency_14 <= sortedFrequencyTemp_13;
      end
    end else if (_T_50) begin
      if (_T_22) begin
        sortedFrequency_14 <= sortedFrequencyTemp_13;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_15 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_23) begin
        sortedFrequency_15 <= sortedFrequencyTemp_14;
      end
    end else if (_T_50) begin
      if (_T_23) begin
        sortedFrequency_15 <= sortedFrequencyTemp_14;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_16 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_24) begin
        sortedFrequency_16 <= sortedFrequencyTemp_15;
      end
    end else if (_T_50) begin
      if (_T_24) begin
        sortedFrequency_16 <= sortedFrequencyTemp_15;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_17 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_25) begin
        sortedFrequency_17 <= sortedFrequencyTemp_16;
      end
    end else if (_T_50) begin
      if (_T_25) begin
        sortedFrequency_17 <= sortedFrequencyTemp_16;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_18 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_26) begin
        sortedFrequency_18 <= sortedFrequencyTemp_17;
      end
    end else if (_T_50) begin
      if (_T_26) begin
        sortedFrequency_18 <= sortedFrequencyTemp_17;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_19 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_27) begin
        sortedFrequency_19 <= sortedFrequencyTemp_18;
      end
    end else if (_T_50) begin
      if (_T_27) begin
        sortedFrequency_19 <= sortedFrequencyTemp_18;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_20 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_28) begin
        sortedFrequency_20 <= sortedFrequencyTemp_19;
      end
    end else if (_T_50) begin
      if (_T_28) begin
        sortedFrequency_20 <= sortedFrequencyTemp_19;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_21 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_29) begin
        sortedFrequency_21 <= sortedFrequencyTemp_20;
      end
    end else if (_T_50) begin
      if (_T_29) begin
        sortedFrequency_21 <= sortedFrequencyTemp_20;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_22 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_30) begin
        sortedFrequency_22 <= sortedFrequencyTemp_21;
      end
    end else if (_T_50) begin
      if (_T_30) begin
        sortedFrequency_22 <= sortedFrequencyTemp_21;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_23 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_31) begin
        sortedFrequency_23 <= sortedFrequencyTemp_22;
      end
    end else if (_T_50) begin
      if (_T_31) begin
        sortedFrequency_23 <= sortedFrequencyTemp_22;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_24 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_32) begin
        sortedFrequency_24 <= sortedFrequencyTemp_23;
      end
    end else if (_T_50) begin
      if (_T_32) begin
        sortedFrequency_24 <= sortedFrequencyTemp_23;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_25 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_33) begin
        sortedFrequency_25 <= sortedFrequencyTemp_24;
      end
    end else if (_T_50) begin
      if (_T_33) begin
        sortedFrequency_25 <= sortedFrequencyTemp_24;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_26 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_34) begin
        sortedFrequency_26 <= sortedFrequencyTemp_25;
      end
    end else if (_T_50) begin
      if (_T_34) begin
        sortedFrequency_26 <= sortedFrequencyTemp_25;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_27 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_35) begin
        sortedFrequency_27 <= sortedFrequencyTemp_26;
      end
    end else if (_T_50) begin
      if (_T_35) begin
        sortedFrequency_27 <= sortedFrequencyTemp_26;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_28 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_36) begin
        sortedFrequency_28 <= sortedFrequencyTemp_27;
      end
    end else if (_T_50) begin
      if (_T_36) begin
        sortedFrequency_28 <= sortedFrequencyTemp_27;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_29 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_37) begin
        sortedFrequency_29 <= sortedFrequencyTemp_28;
      end
    end else if (_T_50) begin
      if (_T_37) begin
        sortedFrequency_29 <= sortedFrequencyTemp_28;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_30 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_38) begin
        sortedFrequency_30 <= sortedFrequencyTemp_29;
      end
    end else if (_T_50) begin
      if (_T_38) begin
        sortedFrequency_30 <= sortedFrequencyTemp_29;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequency_31 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_39) begin
        sortedFrequency_31 <= sortedFrequencyTemp_30;
      end
    end else if (_T_50) begin
      if (_T_39) begin
        sortedFrequency_31 <= sortedFrequencyTemp_30;
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_8) begin
          if (_T) begin
            sortedCharacter_0 <= 9'h0;
          end else if (_T_4) begin
            if (_T_6) begin
              sortedCharacter_0 <= iteration;
            end else begin
              sortedCharacter_0 <= 9'h0;
            end
          end else if (_T_50) begin
            if (_T_51) begin
              sortedCharacter_0 <= 9'h100;
            end else begin
              sortedCharacter_0 <= 9'h0;
            end
          end else begin
            sortedCharacter_0 <= 9'h0;
          end
        end
      end else if (_T_50) begin
        if (_T_8) begin
          if (_T) begin
            sortedCharacter_0 <= 9'h0;
          end else if (_T_4) begin
            if (_T_6) begin
              sortedCharacter_0 <= iteration;
            end else begin
              sortedCharacter_0 <= 9'h0;
            end
          end else if (_T_50) begin
            if (_T_51) begin
              sortedCharacter_0 <= 9'h100;
            end else begin
              sortedCharacter_0 <= 9'h0;
            end
          end else begin
            sortedCharacter_0 <= 9'h0;
          end
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_9) begin
          sortedCharacter_1 <= sortedCharacterTemp_0;
        end
      end else if (_T_50) begin
        if (_T_9) begin
          sortedCharacter_1 <= sortedCharacterTemp_0;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_10) begin
          sortedCharacter_2 <= sortedCharacterTemp_1;
        end
      end else if (_T_50) begin
        if (_T_10) begin
          sortedCharacter_2 <= sortedCharacterTemp_1;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_11) begin
          sortedCharacter_3 <= sortedCharacterTemp_2;
        end
      end else if (_T_50) begin
        if (_T_11) begin
          sortedCharacter_3 <= sortedCharacterTemp_2;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_12) begin
          sortedCharacter_4 <= sortedCharacterTemp_3;
        end
      end else if (_T_50) begin
        if (_T_12) begin
          sortedCharacter_4 <= sortedCharacterTemp_3;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_13) begin
          sortedCharacter_5 <= sortedCharacterTemp_4;
        end
      end else if (_T_50) begin
        if (_T_13) begin
          sortedCharacter_5 <= sortedCharacterTemp_4;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_14) begin
          sortedCharacter_6 <= sortedCharacterTemp_5;
        end
      end else if (_T_50) begin
        if (_T_14) begin
          sortedCharacter_6 <= sortedCharacterTemp_5;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_15) begin
          sortedCharacter_7 <= sortedCharacterTemp_6;
        end
      end else if (_T_50) begin
        if (_T_15) begin
          sortedCharacter_7 <= sortedCharacterTemp_6;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_16) begin
          sortedCharacter_8 <= sortedCharacterTemp_7;
        end
      end else if (_T_50) begin
        if (_T_16) begin
          sortedCharacter_8 <= sortedCharacterTemp_7;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_17) begin
          sortedCharacter_9 <= sortedCharacterTemp_8;
        end
      end else if (_T_50) begin
        if (_T_17) begin
          sortedCharacter_9 <= sortedCharacterTemp_8;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_18) begin
          sortedCharacter_10 <= sortedCharacterTemp_9;
        end
      end else if (_T_50) begin
        if (_T_18) begin
          sortedCharacter_10 <= sortedCharacterTemp_9;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_19) begin
          sortedCharacter_11 <= sortedCharacterTemp_10;
        end
      end else if (_T_50) begin
        if (_T_19) begin
          sortedCharacter_11 <= sortedCharacterTemp_10;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_20) begin
          sortedCharacter_12 <= sortedCharacterTemp_11;
        end
      end else if (_T_50) begin
        if (_T_20) begin
          sortedCharacter_12 <= sortedCharacterTemp_11;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_21) begin
          sortedCharacter_13 <= sortedCharacterTemp_12;
        end
      end else if (_T_50) begin
        if (_T_21) begin
          sortedCharacter_13 <= sortedCharacterTemp_12;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_22) begin
          sortedCharacter_14 <= sortedCharacterTemp_13;
        end
      end else if (_T_50) begin
        if (_T_22) begin
          sortedCharacter_14 <= sortedCharacterTemp_13;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_23) begin
          sortedCharacter_15 <= sortedCharacterTemp_14;
        end
      end else if (_T_50) begin
        if (_T_23) begin
          sortedCharacter_15 <= sortedCharacterTemp_14;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_24) begin
          sortedCharacter_16 <= sortedCharacterTemp_15;
        end
      end else if (_T_50) begin
        if (_T_24) begin
          sortedCharacter_16 <= sortedCharacterTemp_15;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_25) begin
          sortedCharacter_17 <= sortedCharacterTemp_16;
        end
      end else if (_T_50) begin
        if (_T_25) begin
          sortedCharacter_17 <= sortedCharacterTemp_16;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_26) begin
          sortedCharacter_18 <= sortedCharacterTemp_17;
        end
      end else if (_T_50) begin
        if (_T_26) begin
          sortedCharacter_18 <= sortedCharacterTemp_17;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_27) begin
          sortedCharacter_19 <= sortedCharacterTemp_18;
        end
      end else if (_T_50) begin
        if (_T_27) begin
          sortedCharacter_19 <= sortedCharacterTemp_18;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_28) begin
          sortedCharacter_20 <= sortedCharacterTemp_19;
        end
      end else if (_T_50) begin
        if (_T_28) begin
          sortedCharacter_20 <= sortedCharacterTemp_19;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_29) begin
          sortedCharacter_21 <= sortedCharacterTemp_20;
        end
      end else if (_T_50) begin
        if (_T_29) begin
          sortedCharacter_21 <= sortedCharacterTemp_20;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_30) begin
          sortedCharacter_22 <= sortedCharacterTemp_21;
        end
      end else if (_T_50) begin
        if (_T_30) begin
          sortedCharacter_22 <= sortedCharacterTemp_21;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_31) begin
          sortedCharacter_23 <= sortedCharacterTemp_22;
        end
      end else if (_T_50) begin
        if (_T_31) begin
          sortedCharacter_23 <= sortedCharacterTemp_22;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_32) begin
          sortedCharacter_24 <= sortedCharacterTemp_23;
        end
      end else if (_T_50) begin
        if (_T_32) begin
          sortedCharacter_24 <= sortedCharacterTemp_23;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_33) begin
          sortedCharacter_25 <= sortedCharacterTemp_24;
        end
      end else if (_T_50) begin
        if (_T_33) begin
          sortedCharacter_25 <= sortedCharacterTemp_24;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_34) begin
          sortedCharacter_26 <= sortedCharacterTemp_25;
        end
      end else if (_T_50) begin
        if (_T_34) begin
          sortedCharacter_26 <= sortedCharacterTemp_25;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_35) begin
          sortedCharacter_27 <= sortedCharacterTemp_26;
        end
      end else if (_T_50) begin
        if (_T_35) begin
          sortedCharacter_27 <= sortedCharacterTemp_26;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_36) begin
          sortedCharacter_28 <= sortedCharacterTemp_27;
        end
      end else if (_T_50) begin
        if (_T_36) begin
          sortedCharacter_28 <= sortedCharacterTemp_27;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_37) begin
          sortedCharacter_29 <= sortedCharacterTemp_28;
        end
      end else if (_T_50) begin
        if (_T_37) begin
          sortedCharacter_29 <= sortedCharacterTemp_28;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_38) begin
          sortedCharacter_30 <= sortedCharacterTemp_29;
        end
      end else if (_T_50) begin
        if (_T_38) begin
          sortedCharacter_30 <= sortedCharacterTemp_29;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_39) begin
          sortedCharacter_31 <= sortedCharacterTemp_30;
        end
      end else if (_T_50) begin
        if (_T_39) begin
          sortedCharacter_31 <= sortedCharacterTemp_30;
        end
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_0 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_8) begin
        sortedFrequencyTemp_0 <= sortedFrequency_0;
      end else if (_T) begin
        sortedFrequencyTemp_0 <= 13'h0;
      end else if (_T_4) begin
        if (_T_6) begin
          if (8'hff == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_255;
          end else if (8'hfe == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_254;
          end else if (8'hfd == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_253;
          end else if (8'hfc == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_252;
          end else if (8'hfb == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_251;
          end else if (8'hfa == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_250;
          end else if (8'hf9 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_249;
          end else if (8'hf8 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_248;
          end else if (8'hf7 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_247;
          end else if (8'hf6 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_246;
          end else if (8'hf5 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_245;
          end else if (8'hf4 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_244;
          end else if (8'hf3 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_243;
          end else if (8'hf2 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_242;
          end else if (8'hf1 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_241;
          end else if (8'hf0 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_240;
          end else if (8'hef == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_239;
          end else if (8'hee == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_238;
          end else if (8'hed == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_237;
          end else if (8'hec == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_236;
          end else if (8'heb == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_235;
          end else if (8'hea == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_234;
          end else if (8'he9 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_233;
          end else if (8'he8 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_232;
          end else if (8'he7 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_231;
          end else if (8'he6 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_230;
          end else if (8'he5 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_229;
          end else if (8'he4 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_228;
          end else if (8'he3 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_227;
          end else if (8'he2 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_226;
          end else if (8'he1 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_225;
          end else if (8'he0 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_224;
          end else if (8'hdf == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_223;
          end else if (8'hde == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_222;
          end else if (8'hdd == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_221;
          end else if (8'hdc == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_220;
          end else if (8'hdb == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_219;
          end else if (8'hda == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_218;
          end else if (8'hd9 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_217;
          end else if (8'hd8 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_216;
          end else if (8'hd7 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_215;
          end else if (8'hd6 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_214;
          end else if (8'hd5 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_213;
          end else if (8'hd4 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_212;
          end else if (8'hd3 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_211;
          end else if (8'hd2 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_210;
          end else if (8'hd1 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_209;
          end else if (8'hd0 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_208;
          end else if (8'hcf == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_207;
          end else if (8'hce == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_206;
          end else if (8'hcd == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_205;
          end else if (8'hcc == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_204;
          end else if (8'hcb == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_203;
          end else if (8'hca == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_202;
          end else if (8'hc9 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_201;
          end else if (8'hc8 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_200;
          end else if (8'hc7 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_199;
          end else if (8'hc6 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_198;
          end else if (8'hc5 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_197;
          end else if (8'hc4 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_196;
          end else if (8'hc3 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_195;
          end else if (8'hc2 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_194;
          end else if (8'hc1 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_193;
          end else if (8'hc0 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_192;
          end else if (8'hbf == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_191;
          end else if (8'hbe == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_190;
          end else if (8'hbd == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_189;
          end else if (8'hbc == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_188;
          end else if (8'hbb == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_187;
          end else if (8'hba == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_186;
          end else if (8'hb9 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_185;
          end else if (8'hb8 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_184;
          end else if (8'hb7 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_183;
          end else if (8'hb6 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_182;
          end else if (8'hb5 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_181;
          end else if (8'hb4 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_180;
          end else if (8'hb3 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_179;
          end else if (8'hb2 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_178;
          end else if (8'hb1 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_177;
          end else if (8'hb0 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_176;
          end else if (8'haf == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_175;
          end else if (8'hae == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_174;
          end else if (8'had == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_173;
          end else if (8'hac == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_172;
          end else if (8'hab == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_171;
          end else if (8'haa == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_170;
          end else if (8'ha9 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_169;
          end else if (8'ha8 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_168;
          end else if (8'ha7 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_167;
          end else if (8'ha6 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_166;
          end else if (8'ha5 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_165;
          end else if (8'ha4 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_164;
          end else if (8'ha3 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_163;
          end else if (8'ha2 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_162;
          end else if (8'ha1 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_161;
          end else if (8'ha0 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_160;
          end else if (8'h9f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_159;
          end else if (8'h9e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_158;
          end else if (8'h9d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_157;
          end else if (8'h9c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_156;
          end else if (8'h9b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_155;
          end else if (8'h9a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_154;
          end else if (8'h99 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_153;
          end else if (8'h98 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_152;
          end else if (8'h97 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_151;
          end else if (8'h96 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_150;
          end else if (8'h95 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_149;
          end else if (8'h94 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_148;
          end else if (8'h93 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_147;
          end else if (8'h92 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_146;
          end else if (8'h91 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_145;
          end else if (8'h90 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_144;
          end else if (8'h8f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_143;
          end else if (8'h8e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_142;
          end else if (8'h8d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_141;
          end else if (8'h8c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_140;
          end else if (8'h8b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_139;
          end else if (8'h8a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_138;
          end else if (8'h89 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_137;
          end else if (8'h88 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_136;
          end else if (8'h87 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_135;
          end else if (8'h86 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_134;
          end else if (8'h85 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_133;
          end else if (8'h84 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_132;
          end else if (8'h83 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_131;
          end else if (8'h82 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_130;
          end else if (8'h81 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_129;
          end else if (8'h80 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_128;
          end else if (8'h7f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_127;
          end else if (8'h7e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_126;
          end else if (8'h7d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_125;
          end else if (8'h7c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_124;
          end else if (8'h7b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_123;
          end else if (8'h7a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_122;
          end else if (8'h79 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_121;
          end else if (8'h78 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_120;
          end else if (8'h77 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_119;
          end else if (8'h76 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_118;
          end else if (8'h75 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_117;
          end else if (8'h74 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_116;
          end else if (8'h73 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_115;
          end else if (8'h72 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_114;
          end else if (8'h71 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_113;
          end else if (8'h70 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_112;
          end else if (8'h6f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_111;
          end else if (8'h6e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_110;
          end else if (8'h6d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_109;
          end else if (8'h6c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_108;
          end else if (8'h6b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_107;
          end else if (8'h6a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_106;
          end else if (8'h69 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_105;
          end else if (8'h68 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_104;
          end else if (8'h67 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_103;
          end else if (8'h66 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_102;
          end else if (8'h65 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_101;
          end else if (8'h64 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_100;
          end else if (8'h63 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_99;
          end else if (8'h62 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_98;
          end else if (8'h61 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_97;
          end else if (8'h60 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_96;
          end else if (8'h5f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_95;
          end else if (8'h5e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_94;
          end else if (8'h5d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_93;
          end else if (8'h5c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_92;
          end else if (8'h5b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_91;
          end else if (8'h5a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_90;
          end else if (8'h59 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_89;
          end else if (8'h58 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_88;
          end else if (8'h57 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_87;
          end else if (8'h56 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_86;
          end else if (8'h55 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_85;
          end else if (8'h54 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_84;
          end else if (8'h53 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_83;
          end else if (8'h52 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_82;
          end else if (8'h51 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_81;
          end else if (8'h50 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_80;
          end else if (8'h4f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_79;
          end else if (8'h4e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_78;
          end else if (8'h4d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_77;
          end else if (8'h4c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_76;
          end else if (8'h4b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_75;
          end else if (8'h4a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_74;
          end else if (8'h49 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_73;
          end else if (8'h48 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_72;
          end else if (8'h47 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_71;
          end else if (8'h46 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_70;
          end else if (8'h45 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_69;
          end else if (8'h44 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_68;
          end else if (8'h43 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_67;
          end else if (8'h42 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_66;
          end else if (8'h41 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_65;
          end else if (8'h40 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_64;
          end else if (8'h3f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_63;
          end else if (8'h3e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_62;
          end else if (8'h3d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_61;
          end else if (8'h3c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_60;
          end else if (8'h3b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_59;
          end else if (8'h3a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_58;
          end else if (8'h39 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_57;
          end else if (8'h38 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_56;
          end else if (8'h37 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_55;
          end else if (8'h36 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_54;
          end else if (8'h35 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_53;
          end else if (8'h34 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_52;
          end else if (8'h33 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_51;
          end else if (8'h32 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_50;
          end else if (8'h31 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_49;
          end else if (8'h30 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_48;
          end else if (8'h2f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_47;
          end else if (8'h2e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_46;
          end else if (8'h2d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_45;
          end else if (8'h2c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_44;
          end else if (8'h2b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_43;
          end else if (8'h2a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_42;
          end else if (8'h29 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_41;
          end else if (8'h28 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_40;
          end else if (8'h27 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_39;
          end else if (8'h26 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_38;
          end else if (8'h25 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_37;
          end else if (8'h24 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_36;
          end else if (8'h23 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_35;
          end else if (8'h22 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_34;
          end else if (8'h21 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_33;
          end else if (8'h20 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_32;
          end else if (8'h1f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_31;
          end else if (8'h1e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_30;
          end else if (8'h1d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_29;
          end else if (8'h1c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_28;
          end else if (8'h1b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_27;
          end else if (8'h1a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_26;
          end else if (8'h19 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_25;
          end else if (8'h18 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_24;
          end else if (8'h17 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_23;
          end else if (8'h16 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_22;
          end else if (8'h15 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_21;
          end else if (8'h14 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_20;
          end else if (8'h13 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_19;
          end else if (8'h12 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_18;
          end else if (8'h11 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_17;
          end else if (8'h10 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_16;
          end else if (8'hf == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_15;
          end else if (8'he == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_14;
          end else if (8'hd == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_13;
          end else if (8'hc == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_12;
          end else if (8'hb == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_11;
          end else if (8'ha == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_10;
          end else if (8'h9 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_9;
          end else if (8'h8 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_8;
          end else if (8'h7 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_7;
          end else if (8'h6 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_6;
          end else if (8'h5 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_5;
          end else if (8'h4 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_4;
          end else if (8'h3 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_3;
          end else if (8'h2 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_2;
          end else if (8'h1 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_1;
          end else begin
            sortedFrequencyTemp_0 <= io_dataIn_0;
          end
        end else begin
          sortedFrequencyTemp_0 <= 13'h0;
        end
      end else if (_T_50) begin
        if (_T_51) begin
          sortedFrequencyTemp_0 <= escapeFrequency;
        end else begin
          sortedFrequencyTemp_0 <= 13'h0;
        end
      end else begin
        sortedFrequencyTemp_0 <= 13'h0;
      end
    end else if (_T_50) begin
      if (_T_8) begin
        sortedFrequencyTemp_0 <= sortedFrequency_0;
      end else if (_T) begin
        sortedFrequencyTemp_0 <= 13'h0;
      end else if (_T_4) begin
        if (_T_6) begin
          if (8'hff == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_255;
          end else if (8'hfe == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_254;
          end else if (8'hfd == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_253;
          end else if (8'hfc == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_252;
          end else if (8'hfb == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_251;
          end else if (8'hfa == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_250;
          end else if (8'hf9 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_249;
          end else if (8'hf8 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_248;
          end else if (8'hf7 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_247;
          end else if (8'hf6 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_246;
          end else if (8'hf5 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_245;
          end else if (8'hf4 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_244;
          end else if (8'hf3 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_243;
          end else if (8'hf2 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_242;
          end else if (8'hf1 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_241;
          end else if (8'hf0 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_240;
          end else if (8'hef == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_239;
          end else if (8'hee == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_238;
          end else if (8'hed == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_237;
          end else if (8'hec == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_236;
          end else if (8'heb == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_235;
          end else if (8'hea == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_234;
          end else if (8'he9 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_233;
          end else if (8'he8 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_232;
          end else if (8'he7 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_231;
          end else if (8'he6 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_230;
          end else if (8'he5 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_229;
          end else if (8'he4 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_228;
          end else if (8'he3 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_227;
          end else if (8'he2 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_226;
          end else if (8'he1 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_225;
          end else if (8'he0 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_224;
          end else if (8'hdf == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_223;
          end else if (8'hde == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_222;
          end else if (8'hdd == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_221;
          end else if (8'hdc == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_220;
          end else if (8'hdb == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_219;
          end else if (8'hda == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_218;
          end else if (8'hd9 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_217;
          end else if (8'hd8 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_216;
          end else if (8'hd7 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_215;
          end else if (8'hd6 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_214;
          end else if (8'hd5 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_213;
          end else if (8'hd4 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_212;
          end else if (8'hd3 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_211;
          end else if (8'hd2 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_210;
          end else if (8'hd1 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_209;
          end else if (8'hd0 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_208;
          end else if (8'hcf == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_207;
          end else if (8'hce == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_206;
          end else if (8'hcd == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_205;
          end else if (8'hcc == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_204;
          end else if (8'hcb == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_203;
          end else if (8'hca == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_202;
          end else if (8'hc9 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_201;
          end else if (8'hc8 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_200;
          end else if (8'hc7 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_199;
          end else if (8'hc6 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_198;
          end else if (8'hc5 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_197;
          end else if (8'hc4 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_196;
          end else if (8'hc3 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_195;
          end else if (8'hc2 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_194;
          end else if (8'hc1 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_193;
          end else if (8'hc0 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_192;
          end else if (8'hbf == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_191;
          end else if (8'hbe == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_190;
          end else if (8'hbd == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_189;
          end else if (8'hbc == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_188;
          end else if (8'hbb == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_187;
          end else if (8'hba == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_186;
          end else if (8'hb9 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_185;
          end else if (8'hb8 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_184;
          end else if (8'hb7 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_183;
          end else if (8'hb6 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_182;
          end else if (8'hb5 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_181;
          end else if (8'hb4 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_180;
          end else if (8'hb3 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_179;
          end else if (8'hb2 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_178;
          end else if (8'hb1 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_177;
          end else if (8'hb0 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_176;
          end else if (8'haf == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_175;
          end else if (8'hae == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_174;
          end else if (8'had == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_173;
          end else if (8'hac == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_172;
          end else if (8'hab == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_171;
          end else if (8'haa == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_170;
          end else if (8'ha9 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_169;
          end else if (8'ha8 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_168;
          end else if (8'ha7 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_167;
          end else if (8'ha6 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_166;
          end else if (8'ha5 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_165;
          end else if (8'ha4 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_164;
          end else if (8'ha3 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_163;
          end else if (8'ha2 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_162;
          end else if (8'ha1 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_161;
          end else if (8'ha0 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_160;
          end else if (8'h9f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_159;
          end else if (8'h9e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_158;
          end else if (8'h9d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_157;
          end else if (8'h9c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_156;
          end else if (8'h9b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_155;
          end else if (8'h9a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_154;
          end else if (8'h99 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_153;
          end else if (8'h98 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_152;
          end else if (8'h97 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_151;
          end else if (8'h96 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_150;
          end else if (8'h95 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_149;
          end else if (8'h94 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_148;
          end else if (8'h93 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_147;
          end else if (8'h92 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_146;
          end else if (8'h91 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_145;
          end else if (8'h90 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_144;
          end else if (8'h8f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_143;
          end else if (8'h8e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_142;
          end else if (8'h8d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_141;
          end else if (8'h8c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_140;
          end else if (8'h8b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_139;
          end else if (8'h8a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_138;
          end else if (8'h89 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_137;
          end else if (8'h88 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_136;
          end else if (8'h87 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_135;
          end else if (8'h86 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_134;
          end else if (8'h85 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_133;
          end else if (8'h84 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_132;
          end else if (8'h83 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_131;
          end else if (8'h82 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_130;
          end else if (8'h81 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_129;
          end else if (8'h80 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_128;
          end else if (8'h7f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_127;
          end else if (8'h7e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_126;
          end else if (8'h7d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_125;
          end else if (8'h7c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_124;
          end else if (8'h7b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_123;
          end else if (8'h7a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_122;
          end else if (8'h79 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_121;
          end else if (8'h78 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_120;
          end else if (8'h77 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_119;
          end else if (8'h76 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_118;
          end else if (8'h75 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_117;
          end else if (8'h74 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_116;
          end else if (8'h73 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_115;
          end else if (8'h72 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_114;
          end else if (8'h71 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_113;
          end else if (8'h70 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_112;
          end else if (8'h6f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_111;
          end else if (8'h6e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_110;
          end else if (8'h6d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_109;
          end else if (8'h6c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_108;
          end else if (8'h6b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_107;
          end else if (8'h6a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_106;
          end else if (8'h69 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_105;
          end else if (8'h68 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_104;
          end else if (8'h67 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_103;
          end else if (8'h66 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_102;
          end else if (8'h65 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_101;
          end else if (8'h64 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_100;
          end else if (8'h63 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_99;
          end else if (8'h62 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_98;
          end else if (8'h61 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_97;
          end else if (8'h60 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_96;
          end else if (8'h5f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_95;
          end else if (8'h5e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_94;
          end else if (8'h5d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_93;
          end else if (8'h5c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_92;
          end else if (8'h5b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_91;
          end else if (8'h5a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_90;
          end else if (8'h59 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_89;
          end else if (8'h58 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_88;
          end else if (8'h57 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_87;
          end else if (8'h56 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_86;
          end else if (8'h55 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_85;
          end else if (8'h54 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_84;
          end else if (8'h53 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_83;
          end else if (8'h52 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_82;
          end else if (8'h51 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_81;
          end else if (8'h50 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_80;
          end else if (8'h4f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_79;
          end else if (8'h4e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_78;
          end else if (8'h4d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_77;
          end else if (8'h4c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_76;
          end else if (8'h4b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_75;
          end else if (8'h4a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_74;
          end else if (8'h49 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_73;
          end else if (8'h48 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_72;
          end else if (8'h47 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_71;
          end else if (8'h46 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_70;
          end else if (8'h45 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_69;
          end else if (8'h44 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_68;
          end else if (8'h43 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_67;
          end else if (8'h42 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_66;
          end else if (8'h41 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_65;
          end else if (8'h40 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_64;
          end else if (8'h3f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_63;
          end else if (8'h3e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_62;
          end else if (8'h3d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_61;
          end else if (8'h3c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_60;
          end else if (8'h3b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_59;
          end else if (8'h3a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_58;
          end else if (8'h39 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_57;
          end else if (8'h38 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_56;
          end else if (8'h37 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_55;
          end else if (8'h36 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_54;
          end else if (8'h35 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_53;
          end else if (8'h34 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_52;
          end else if (8'h33 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_51;
          end else if (8'h32 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_50;
          end else if (8'h31 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_49;
          end else if (8'h30 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_48;
          end else if (8'h2f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_47;
          end else if (8'h2e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_46;
          end else if (8'h2d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_45;
          end else if (8'h2c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_44;
          end else if (8'h2b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_43;
          end else if (8'h2a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_42;
          end else if (8'h29 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_41;
          end else if (8'h28 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_40;
          end else if (8'h27 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_39;
          end else if (8'h26 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_38;
          end else if (8'h25 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_37;
          end else if (8'h24 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_36;
          end else if (8'h23 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_35;
          end else if (8'h22 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_34;
          end else if (8'h21 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_33;
          end else if (8'h20 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_32;
          end else if (8'h1f == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_31;
          end else if (8'h1e == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_30;
          end else if (8'h1d == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_29;
          end else if (8'h1c == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_28;
          end else if (8'h1b == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_27;
          end else if (8'h1a == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_26;
          end else if (8'h19 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_25;
          end else if (8'h18 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_24;
          end else if (8'h17 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_23;
          end else if (8'h16 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_22;
          end else if (8'h15 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_21;
          end else if (8'h14 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_20;
          end else if (8'h13 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_19;
          end else if (8'h12 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_18;
          end else if (8'h11 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_17;
          end else if (8'h10 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_16;
          end else if (8'hf == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_15;
          end else if (8'he == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_14;
          end else if (8'hd == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_13;
          end else if (8'hc == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_12;
          end else if (8'hb == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_11;
          end else if (8'ha == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_10;
          end else if (8'h9 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_9;
          end else if (8'h8 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_8;
          end else if (8'h7 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_7;
          end else if (8'h6 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_6;
          end else if (8'h5 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_5;
          end else if (8'h4 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_4;
          end else if (8'h3 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_3;
          end else if (8'h2 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_2;
          end else if (8'h1 == iteration[7:0]) begin
            sortedFrequencyTemp_0 <= io_dataIn_1;
          end else begin
            sortedFrequencyTemp_0 <= io_dataIn_0;
          end
        end else begin
          sortedFrequencyTemp_0 <= 13'h0;
        end
      end else if (_T_50) begin
        if (_T_51) begin
          sortedFrequencyTemp_0 <= escapeFrequency;
        end else begin
          sortedFrequencyTemp_0 <= 13'h0;
        end
      end else begin
        sortedFrequencyTemp_0 <= 13'h0;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_1 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_9) begin
        sortedFrequencyTemp_1 <= sortedFrequency_1;
      end else begin
        sortedFrequencyTemp_1 <= sortedFrequencyTemp_0;
      end
    end else if (_T_50) begin
      if (_T_9) begin
        sortedFrequencyTemp_1 <= sortedFrequency_1;
      end else begin
        sortedFrequencyTemp_1 <= sortedFrequencyTemp_0;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_2 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_10) begin
        sortedFrequencyTemp_2 <= sortedFrequency_2;
      end else begin
        sortedFrequencyTemp_2 <= sortedFrequencyTemp_1;
      end
    end else if (_T_50) begin
      if (_T_10) begin
        sortedFrequencyTemp_2 <= sortedFrequency_2;
      end else begin
        sortedFrequencyTemp_2 <= sortedFrequencyTemp_1;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_3 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_11) begin
        sortedFrequencyTemp_3 <= sortedFrequency_3;
      end else begin
        sortedFrequencyTemp_3 <= sortedFrequencyTemp_2;
      end
    end else if (_T_50) begin
      if (_T_11) begin
        sortedFrequencyTemp_3 <= sortedFrequency_3;
      end else begin
        sortedFrequencyTemp_3 <= sortedFrequencyTemp_2;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_4 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_12) begin
        sortedFrequencyTemp_4 <= sortedFrequency_4;
      end else begin
        sortedFrequencyTemp_4 <= sortedFrequencyTemp_3;
      end
    end else if (_T_50) begin
      if (_T_12) begin
        sortedFrequencyTemp_4 <= sortedFrequency_4;
      end else begin
        sortedFrequencyTemp_4 <= sortedFrequencyTemp_3;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_5 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_13) begin
        sortedFrequencyTemp_5 <= sortedFrequency_5;
      end else begin
        sortedFrequencyTemp_5 <= sortedFrequencyTemp_4;
      end
    end else if (_T_50) begin
      if (_T_13) begin
        sortedFrequencyTemp_5 <= sortedFrequency_5;
      end else begin
        sortedFrequencyTemp_5 <= sortedFrequencyTemp_4;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_6 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_14) begin
        sortedFrequencyTemp_6 <= sortedFrequency_6;
      end else begin
        sortedFrequencyTemp_6 <= sortedFrequencyTemp_5;
      end
    end else if (_T_50) begin
      if (_T_14) begin
        sortedFrequencyTemp_6 <= sortedFrequency_6;
      end else begin
        sortedFrequencyTemp_6 <= sortedFrequencyTemp_5;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_7 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_15) begin
        sortedFrequencyTemp_7 <= sortedFrequency_7;
      end else begin
        sortedFrequencyTemp_7 <= sortedFrequencyTemp_6;
      end
    end else if (_T_50) begin
      if (_T_15) begin
        sortedFrequencyTemp_7 <= sortedFrequency_7;
      end else begin
        sortedFrequencyTemp_7 <= sortedFrequencyTemp_6;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_8 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_16) begin
        sortedFrequencyTemp_8 <= sortedFrequency_8;
      end else begin
        sortedFrequencyTemp_8 <= sortedFrequencyTemp_7;
      end
    end else if (_T_50) begin
      if (_T_16) begin
        sortedFrequencyTemp_8 <= sortedFrequency_8;
      end else begin
        sortedFrequencyTemp_8 <= sortedFrequencyTemp_7;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_9 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_17) begin
        sortedFrequencyTemp_9 <= sortedFrequency_9;
      end else begin
        sortedFrequencyTemp_9 <= sortedFrequencyTemp_8;
      end
    end else if (_T_50) begin
      if (_T_17) begin
        sortedFrequencyTemp_9 <= sortedFrequency_9;
      end else begin
        sortedFrequencyTemp_9 <= sortedFrequencyTemp_8;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_10 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_18) begin
        sortedFrequencyTemp_10 <= sortedFrequency_10;
      end else begin
        sortedFrequencyTemp_10 <= sortedFrequencyTemp_9;
      end
    end else if (_T_50) begin
      if (_T_18) begin
        sortedFrequencyTemp_10 <= sortedFrequency_10;
      end else begin
        sortedFrequencyTemp_10 <= sortedFrequencyTemp_9;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_11 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_19) begin
        sortedFrequencyTemp_11 <= sortedFrequency_11;
      end else begin
        sortedFrequencyTemp_11 <= sortedFrequencyTemp_10;
      end
    end else if (_T_50) begin
      if (_T_19) begin
        sortedFrequencyTemp_11 <= sortedFrequency_11;
      end else begin
        sortedFrequencyTemp_11 <= sortedFrequencyTemp_10;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_12 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_20) begin
        sortedFrequencyTemp_12 <= sortedFrequency_12;
      end else begin
        sortedFrequencyTemp_12 <= sortedFrequencyTemp_11;
      end
    end else if (_T_50) begin
      if (_T_20) begin
        sortedFrequencyTemp_12 <= sortedFrequency_12;
      end else begin
        sortedFrequencyTemp_12 <= sortedFrequencyTemp_11;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_13 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_21) begin
        sortedFrequencyTemp_13 <= sortedFrequency_13;
      end else begin
        sortedFrequencyTemp_13 <= sortedFrequencyTemp_12;
      end
    end else if (_T_50) begin
      if (_T_21) begin
        sortedFrequencyTemp_13 <= sortedFrequency_13;
      end else begin
        sortedFrequencyTemp_13 <= sortedFrequencyTemp_12;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_14 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_22) begin
        sortedFrequencyTemp_14 <= sortedFrequency_14;
      end else begin
        sortedFrequencyTemp_14 <= sortedFrequencyTemp_13;
      end
    end else if (_T_50) begin
      if (_T_22) begin
        sortedFrequencyTemp_14 <= sortedFrequency_14;
      end else begin
        sortedFrequencyTemp_14 <= sortedFrequencyTemp_13;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_15 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_23) begin
        sortedFrequencyTemp_15 <= sortedFrequency_15;
      end else begin
        sortedFrequencyTemp_15 <= sortedFrequencyTemp_14;
      end
    end else if (_T_50) begin
      if (_T_23) begin
        sortedFrequencyTemp_15 <= sortedFrequency_15;
      end else begin
        sortedFrequencyTemp_15 <= sortedFrequencyTemp_14;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_16 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_24) begin
        sortedFrequencyTemp_16 <= sortedFrequency_16;
      end else begin
        sortedFrequencyTemp_16 <= sortedFrequencyTemp_15;
      end
    end else if (_T_50) begin
      if (_T_24) begin
        sortedFrequencyTemp_16 <= sortedFrequency_16;
      end else begin
        sortedFrequencyTemp_16 <= sortedFrequencyTemp_15;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_17 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_25) begin
        sortedFrequencyTemp_17 <= sortedFrequency_17;
      end else begin
        sortedFrequencyTemp_17 <= sortedFrequencyTemp_16;
      end
    end else if (_T_50) begin
      if (_T_25) begin
        sortedFrequencyTemp_17 <= sortedFrequency_17;
      end else begin
        sortedFrequencyTemp_17 <= sortedFrequencyTemp_16;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_18 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_26) begin
        sortedFrequencyTemp_18 <= sortedFrequency_18;
      end else begin
        sortedFrequencyTemp_18 <= sortedFrequencyTemp_17;
      end
    end else if (_T_50) begin
      if (_T_26) begin
        sortedFrequencyTemp_18 <= sortedFrequency_18;
      end else begin
        sortedFrequencyTemp_18 <= sortedFrequencyTemp_17;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_19 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_27) begin
        sortedFrequencyTemp_19 <= sortedFrequency_19;
      end else begin
        sortedFrequencyTemp_19 <= sortedFrequencyTemp_18;
      end
    end else if (_T_50) begin
      if (_T_27) begin
        sortedFrequencyTemp_19 <= sortedFrequency_19;
      end else begin
        sortedFrequencyTemp_19 <= sortedFrequencyTemp_18;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_20 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_28) begin
        sortedFrequencyTemp_20 <= sortedFrequency_20;
      end else begin
        sortedFrequencyTemp_20 <= sortedFrequencyTemp_19;
      end
    end else if (_T_50) begin
      if (_T_28) begin
        sortedFrequencyTemp_20 <= sortedFrequency_20;
      end else begin
        sortedFrequencyTemp_20 <= sortedFrequencyTemp_19;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_21 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_29) begin
        sortedFrequencyTemp_21 <= sortedFrequency_21;
      end else begin
        sortedFrequencyTemp_21 <= sortedFrequencyTemp_20;
      end
    end else if (_T_50) begin
      if (_T_29) begin
        sortedFrequencyTemp_21 <= sortedFrequency_21;
      end else begin
        sortedFrequencyTemp_21 <= sortedFrequencyTemp_20;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_22 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_30) begin
        sortedFrequencyTemp_22 <= sortedFrequency_22;
      end else begin
        sortedFrequencyTemp_22 <= sortedFrequencyTemp_21;
      end
    end else if (_T_50) begin
      if (_T_30) begin
        sortedFrequencyTemp_22 <= sortedFrequency_22;
      end else begin
        sortedFrequencyTemp_22 <= sortedFrequencyTemp_21;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_23 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_31) begin
        sortedFrequencyTemp_23 <= sortedFrequency_23;
      end else begin
        sortedFrequencyTemp_23 <= sortedFrequencyTemp_22;
      end
    end else if (_T_50) begin
      if (_T_31) begin
        sortedFrequencyTemp_23 <= sortedFrequency_23;
      end else begin
        sortedFrequencyTemp_23 <= sortedFrequencyTemp_22;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_24 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_32) begin
        sortedFrequencyTemp_24 <= sortedFrequency_24;
      end else begin
        sortedFrequencyTemp_24 <= sortedFrequencyTemp_23;
      end
    end else if (_T_50) begin
      if (_T_32) begin
        sortedFrequencyTemp_24 <= sortedFrequency_24;
      end else begin
        sortedFrequencyTemp_24 <= sortedFrequencyTemp_23;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_25 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_33) begin
        sortedFrequencyTemp_25 <= sortedFrequency_25;
      end else begin
        sortedFrequencyTemp_25 <= sortedFrequencyTemp_24;
      end
    end else if (_T_50) begin
      if (_T_33) begin
        sortedFrequencyTemp_25 <= sortedFrequency_25;
      end else begin
        sortedFrequencyTemp_25 <= sortedFrequencyTemp_24;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_26 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_34) begin
        sortedFrequencyTemp_26 <= sortedFrequency_26;
      end else begin
        sortedFrequencyTemp_26 <= sortedFrequencyTemp_25;
      end
    end else if (_T_50) begin
      if (_T_34) begin
        sortedFrequencyTemp_26 <= sortedFrequency_26;
      end else begin
        sortedFrequencyTemp_26 <= sortedFrequencyTemp_25;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_27 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_35) begin
        sortedFrequencyTemp_27 <= sortedFrequency_27;
      end else begin
        sortedFrequencyTemp_27 <= sortedFrequencyTemp_26;
      end
    end else if (_T_50) begin
      if (_T_35) begin
        sortedFrequencyTemp_27 <= sortedFrequency_27;
      end else begin
        sortedFrequencyTemp_27 <= sortedFrequencyTemp_26;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_28 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_36) begin
        sortedFrequencyTemp_28 <= sortedFrequency_28;
      end else begin
        sortedFrequencyTemp_28 <= sortedFrequencyTemp_27;
      end
    end else if (_T_50) begin
      if (_T_36) begin
        sortedFrequencyTemp_28 <= sortedFrequency_28;
      end else begin
        sortedFrequencyTemp_28 <= sortedFrequencyTemp_27;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_29 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_37) begin
        sortedFrequencyTemp_29 <= sortedFrequency_29;
      end else begin
        sortedFrequencyTemp_29 <= sortedFrequencyTemp_28;
      end
    end else if (_T_50) begin
      if (_T_37) begin
        sortedFrequencyTemp_29 <= sortedFrequency_29;
      end else begin
        sortedFrequencyTemp_29 <= sortedFrequencyTemp_28;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedFrequencyTemp_30 <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_38) begin
        sortedFrequencyTemp_30 <= sortedFrequency_30;
      end else begin
        sortedFrequencyTemp_30 <= sortedFrequencyTemp_29;
      end
    end else if (_T_50) begin
      if (_T_38) begin
        sortedFrequencyTemp_30 <= sortedFrequency_30;
      end else begin
        sortedFrequencyTemp_30 <= sortedFrequencyTemp_29;
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_8) begin
          sortedCharacterTemp_0 <= sortedCharacter_0;
        end else if (_T) begin
          sortedCharacterTemp_0 <= 9'h0;
        end else if (_T_4) begin
          if (_T_6) begin
            sortedCharacterTemp_0 <= iteration;
          end else begin
            sortedCharacterTemp_0 <= 9'h0;
          end
        end else if (_T_50) begin
          if (_T_51) begin
            sortedCharacterTemp_0 <= 9'h100;
          end else begin
            sortedCharacterTemp_0 <= 9'h0;
          end
        end else begin
          sortedCharacterTemp_0 <= 9'h0;
        end
      end else if (_T_50) begin
        if (_T_8) begin
          sortedCharacterTemp_0 <= sortedCharacter_0;
        end else if (_T) begin
          sortedCharacterTemp_0 <= 9'h0;
        end else if (_T_4) begin
          if (_T_6) begin
            sortedCharacterTemp_0 <= iteration;
          end else begin
            sortedCharacterTemp_0 <= 9'h0;
          end
        end else if (_T_50) begin
          if (_T_51) begin
            sortedCharacterTemp_0 <= 9'h100;
          end else begin
            sortedCharacterTemp_0 <= 9'h0;
          end
        end else begin
          sortedCharacterTemp_0 <= 9'h0;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_9) begin
          sortedCharacterTemp_1 <= sortedCharacter_1;
        end else begin
          sortedCharacterTemp_1 <= sortedCharacterTemp_0;
        end
      end else if (_T_50) begin
        if (_T_9) begin
          sortedCharacterTemp_1 <= sortedCharacter_1;
        end else begin
          sortedCharacterTemp_1 <= sortedCharacterTemp_0;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_10) begin
          sortedCharacterTemp_2 <= sortedCharacter_2;
        end else begin
          sortedCharacterTemp_2 <= sortedCharacterTemp_1;
        end
      end else if (_T_50) begin
        if (_T_10) begin
          sortedCharacterTemp_2 <= sortedCharacter_2;
        end else begin
          sortedCharacterTemp_2 <= sortedCharacterTemp_1;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_11) begin
          sortedCharacterTemp_3 <= sortedCharacter_3;
        end else begin
          sortedCharacterTemp_3 <= sortedCharacterTemp_2;
        end
      end else if (_T_50) begin
        if (_T_11) begin
          sortedCharacterTemp_3 <= sortedCharacter_3;
        end else begin
          sortedCharacterTemp_3 <= sortedCharacterTemp_2;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_12) begin
          sortedCharacterTemp_4 <= sortedCharacter_4;
        end else begin
          sortedCharacterTemp_4 <= sortedCharacterTemp_3;
        end
      end else if (_T_50) begin
        if (_T_12) begin
          sortedCharacterTemp_4 <= sortedCharacter_4;
        end else begin
          sortedCharacterTemp_4 <= sortedCharacterTemp_3;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_13) begin
          sortedCharacterTemp_5 <= sortedCharacter_5;
        end else begin
          sortedCharacterTemp_5 <= sortedCharacterTemp_4;
        end
      end else if (_T_50) begin
        if (_T_13) begin
          sortedCharacterTemp_5 <= sortedCharacter_5;
        end else begin
          sortedCharacterTemp_5 <= sortedCharacterTemp_4;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_14) begin
          sortedCharacterTemp_6 <= sortedCharacter_6;
        end else begin
          sortedCharacterTemp_6 <= sortedCharacterTemp_5;
        end
      end else if (_T_50) begin
        if (_T_14) begin
          sortedCharacterTemp_6 <= sortedCharacter_6;
        end else begin
          sortedCharacterTemp_6 <= sortedCharacterTemp_5;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_15) begin
          sortedCharacterTemp_7 <= sortedCharacter_7;
        end else begin
          sortedCharacterTemp_7 <= sortedCharacterTemp_6;
        end
      end else if (_T_50) begin
        if (_T_15) begin
          sortedCharacterTemp_7 <= sortedCharacter_7;
        end else begin
          sortedCharacterTemp_7 <= sortedCharacterTemp_6;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_16) begin
          sortedCharacterTemp_8 <= sortedCharacter_8;
        end else begin
          sortedCharacterTemp_8 <= sortedCharacterTemp_7;
        end
      end else if (_T_50) begin
        if (_T_16) begin
          sortedCharacterTemp_8 <= sortedCharacter_8;
        end else begin
          sortedCharacterTemp_8 <= sortedCharacterTemp_7;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_17) begin
          sortedCharacterTemp_9 <= sortedCharacter_9;
        end else begin
          sortedCharacterTemp_9 <= sortedCharacterTemp_8;
        end
      end else if (_T_50) begin
        if (_T_17) begin
          sortedCharacterTemp_9 <= sortedCharacter_9;
        end else begin
          sortedCharacterTemp_9 <= sortedCharacterTemp_8;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_18) begin
          sortedCharacterTemp_10 <= sortedCharacter_10;
        end else begin
          sortedCharacterTemp_10 <= sortedCharacterTemp_9;
        end
      end else if (_T_50) begin
        if (_T_18) begin
          sortedCharacterTemp_10 <= sortedCharacter_10;
        end else begin
          sortedCharacterTemp_10 <= sortedCharacterTemp_9;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_19) begin
          sortedCharacterTemp_11 <= sortedCharacter_11;
        end else begin
          sortedCharacterTemp_11 <= sortedCharacterTemp_10;
        end
      end else if (_T_50) begin
        if (_T_19) begin
          sortedCharacterTemp_11 <= sortedCharacter_11;
        end else begin
          sortedCharacterTemp_11 <= sortedCharacterTemp_10;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_20) begin
          sortedCharacterTemp_12 <= sortedCharacter_12;
        end else begin
          sortedCharacterTemp_12 <= sortedCharacterTemp_11;
        end
      end else if (_T_50) begin
        if (_T_20) begin
          sortedCharacterTemp_12 <= sortedCharacter_12;
        end else begin
          sortedCharacterTemp_12 <= sortedCharacterTemp_11;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_21) begin
          sortedCharacterTemp_13 <= sortedCharacter_13;
        end else begin
          sortedCharacterTemp_13 <= sortedCharacterTemp_12;
        end
      end else if (_T_50) begin
        if (_T_21) begin
          sortedCharacterTemp_13 <= sortedCharacter_13;
        end else begin
          sortedCharacterTemp_13 <= sortedCharacterTemp_12;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_22) begin
          sortedCharacterTemp_14 <= sortedCharacter_14;
        end else begin
          sortedCharacterTemp_14 <= sortedCharacterTemp_13;
        end
      end else if (_T_50) begin
        if (_T_22) begin
          sortedCharacterTemp_14 <= sortedCharacter_14;
        end else begin
          sortedCharacterTemp_14 <= sortedCharacterTemp_13;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_23) begin
          sortedCharacterTemp_15 <= sortedCharacter_15;
        end else begin
          sortedCharacterTemp_15 <= sortedCharacterTemp_14;
        end
      end else if (_T_50) begin
        if (_T_23) begin
          sortedCharacterTemp_15 <= sortedCharacter_15;
        end else begin
          sortedCharacterTemp_15 <= sortedCharacterTemp_14;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_24) begin
          sortedCharacterTemp_16 <= sortedCharacter_16;
        end else begin
          sortedCharacterTemp_16 <= sortedCharacterTemp_15;
        end
      end else if (_T_50) begin
        if (_T_24) begin
          sortedCharacterTemp_16 <= sortedCharacter_16;
        end else begin
          sortedCharacterTemp_16 <= sortedCharacterTemp_15;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_25) begin
          sortedCharacterTemp_17 <= sortedCharacter_17;
        end else begin
          sortedCharacterTemp_17 <= sortedCharacterTemp_16;
        end
      end else if (_T_50) begin
        if (_T_25) begin
          sortedCharacterTemp_17 <= sortedCharacter_17;
        end else begin
          sortedCharacterTemp_17 <= sortedCharacterTemp_16;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_26) begin
          sortedCharacterTemp_18 <= sortedCharacter_18;
        end else begin
          sortedCharacterTemp_18 <= sortedCharacterTemp_17;
        end
      end else if (_T_50) begin
        if (_T_26) begin
          sortedCharacterTemp_18 <= sortedCharacter_18;
        end else begin
          sortedCharacterTemp_18 <= sortedCharacterTemp_17;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_27) begin
          sortedCharacterTemp_19 <= sortedCharacter_19;
        end else begin
          sortedCharacterTemp_19 <= sortedCharacterTemp_18;
        end
      end else if (_T_50) begin
        if (_T_27) begin
          sortedCharacterTemp_19 <= sortedCharacter_19;
        end else begin
          sortedCharacterTemp_19 <= sortedCharacterTemp_18;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_28) begin
          sortedCharacterTemp_20 <= sortedCharacter_20;
        end else begin
          sortedCharacterTemp_20 <= sortedCharacterTemp_19;
        end
      end else if (_T_50) begin
        if (_T_28) begin
          sortedCharacterTemp_20 <= sortedCharacter_20;
        end else begin
          sortedCharacterTemp_20 <= sortedCharacterTemp_19;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_29) begin
          sortedCharacterTemp_21 <= sortedCharacter_21;
        end else begin
          sortedCharacterTemp_21 <= sortedCharacterTemp_20;
        end
      end else if (_T_50) begin
        if (_T_29) begin
          sortedCharacterTemp_21 <= sortedCharacter_21;
        end else begin
          sortedCharacterTemp_21 <= sortedCharacterTemp_20;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_30) begin
          sortedCharacterTemp_22 <= sortedCharacter_22;
        end else begin
          sortedCharacterTemp_22 <= sortedCharacterTemp_21;
        end
      end else if (_T_50) begin
        if (_T_30) begin
          sortedCharacterTemp_22 <= sortedCharacter_22;
        end else begin
          sortedCharacterTemp_22 <= sortedCharacterTemp_21;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_31) begin
          sortedCharacterTemp_23 <= sortedCharacter_23;
        end else begin
          sortedCharacterTemp_23 <= sortedCharacterTemp_22;
        end
      end else if (_T_50) begin
        if (_T_31) begin
          sortedCharacterTemp_23 <= sortedCharacter_23;
        end else begin
          sortedCharacterTemp_23 <= sortedCharacterTemp_22;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_32) begin
          sortedCharacterTemp_24 <= sortedCharacter_24;
        end else begin
          sortedCharacterTemp_24 <= sortedCharacterTemp_23;
        end
      end else if (_T_50) begin
        if (_T_32) begin
          sortedCharacterTemp_24 <= sortedCharacter_24;
        end else begin
          sortedCharacterTemp_24 <= sortedCharacterTemp_23;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_33) begin
          sortedCharacterTemp_25 <= sortedCharacter_25;
        end else begin
          sortedCharacterTemp_25 <= sortedCharacterTemp_24;
        end
      end else if (_T_50) begin
        if (_T_33) begin
          sortedCharacterTemp_25 <= sortedCharacter_25;
        end else begin
          sortedCharacterTemp_25 <= sortedCharacterTemp_24;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_34) begin
          sortedCharacterTemp_26 <= sortedCharacter_26;
        end else begin
          sortedCharacterTemp_26 <= sortedCharacterTemp_25;
        end
      end else if (_T_50) begin
        if (_T_34) begin
          sortedCharacterTemp_26 <= sortedCharacter_26;
        end else begin
          sortedCharacterTemp_26 <= sortedCharacterTemp_25;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_35) begin
          sortedCharacterTemp_27 <= sortedCharacter_27;
        end else begin
          sortedCharacterTemp_27 <= sortedCharacterTemp_26;
        end
      end else if (_T_50) begin
        if (_T_35) begin
          sortedCharacterTemp_27 <= sortedCharacter_27;
        end else begin
          sortedCharacterTemp_27 <= sortedCharacterTemp_26;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_36) begin
          sortedCharacterTemp_28 <= sortedCharacter_28;
        end else begin
          sortedCharacterTemp_28 <= sortedCharacterTemp_27;
        end
      end else if (_T_50) begin
        if (_T_36) begin
          sortedCharacterTemp_28 <= sortedCharacter_28;
        end else begin
          sortedCharacterTemp_28 <= sortedCharacterTemp_27;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_37) begin
          sortedCharacterTemp_29 <= sortedCharacter_29;
        end else begin
          sortedCharacterTemp_29 <= sortedCharacterTemp_28;
        end
      end else if (_T_50) begin
        if (_T_37) begin
          sortedCharacterTemp_29 <= sortedCharacter_29;
        end else begin
          sortedCharacterTemp_29 <= sortedCharacterTemp_28;
        end
      end
    end
    if (!(_T)) begin
      if (_T_4) begin
        if (_T_38) begin
          sortedCharacterTemp_30 <= sortedCharacter_30;
        end else begin
          sortedCharacterTemp_30 <= sortedCharacterTemp_29;
        end
      end else if (_T_50) begin
        if (_T_38) begin
          sortedCharacterTemp_30 <= sortedCharacter_30;
        end else begin
          sortedCharacterTemp_30 <= sortedCharacterTemp_29;
        end
      end
    end
    if (_T) begin
      if (io_start) begin
        escapeFrequency <= 13'h0;
      end
    end else if (_T_4) begin
      if (_T_46) begin
        if (_T_47) begin
          escapeFrequency <= _T_41;
        end else if (_T_39) begin
          escapeFrequency <= _T_41;
        end else begin
          escapeFrequency <= _T_43;
        end
      end else if (_T_39) begin
        escapeFrequency <= _T_41;
      end else begin
        escapeFrequency <= _T_43;
      end
    end
  end
endmodule
module characterFrequencyModule(
  input         clock,
  input         reset,
  input         io_start,
  output [11:0] io_input_currentByteOut,
  input  [7:0]  io_input_dataIn_0,
  input         io_input_valid,
  output        io_input_ready,
  output [12:0] io_outputs_sortedFrequency_0,
  output [12:0] io_outputs_sortedFrequency_1,
  output [12:0] io_outputs_sortedFrequency_2,
  output [12:0] io_outputs_sortedFrequency_3,
  output [12:0] io_outputs_sortedFrequency_4,
  output [12:0] io_outputs_sortedFrequency_5,
  output [12:0] io_outputs_sortedFrequency_6,
  output [12:0] io_outputs_sortedFrequency_7,
  output [12:0] io_outputs_sortedFrequency_8,
  output [12:0] io_outputs_sortedFrequency_9,
  output [12:0] io_outputs_sortedFrequency_10,
  output [12:0] io_outputs_sortedFrequency_11,
  output [12:0] io_outputs_sortedFrequency_12,
  output [12:0] io_outputs_sortedFrequency_13,
  output [12:0] io_outputs_sortedFrequency_14,
  output [12:0] io_outputs_sortedFrequency_15,
  output [12:0] io_outputs_sortedFrequency_16,
  output [12:0] io_outputs_sortedFrequency_17,
  output [12:0] io_outputs_sortedFrequency_18,
  output [12:0] io_outputs_sortedFrequency_19,
  output [12:0] io_outputs_sortedFrequency_20,
  output [12:0] io_outputs_sortedFrequency_21,
  output [12:0] io_outputs_sortedFrequency_22,
  output [12:0] io_outputs_sortedFrequency_23,
  output [12:0] io_outputs_sortedFrequency_24,
  output [12:0] io_outputs_sortedFrequency_25,
  output [12:0] io_outputs_sortedFrequency_26,
  output [12:0] io_outputs_sortedFrequency_27,
  output [12:0] io_outputs_sortedFrequency_28,
  output [12:0] io_outputs_sortedFrequency_29,
  output [12:0] io_outputs_sortedFrequency_30,
  output [12:0] io_outputs_sortedFrequency_31,
  output [8:0]  io_outputs_sortedCharacter_0,
  output [8:0]  io_outputs_sortedCharacter_1,
  output [8:0]  io_outputs_sortedCharacter_2,
  output [8:0]  io_outputs_sortedCharacter_3,
  output [8:0]  io_outputs_sortedCharacter_4,
  output [8:0]  io_outputs_sortedCharacter_5,
  output [8:0]  io_outputs_sortedCharacter_6,
  output [8:0]  io_outputs_sortedCharacter_7,
  output [8:0]  io_outputs_sortedCharacter_8,
  output [8:0]  io_outputs_sortedCharacter_9,
  output [8:0]  io_outputs_sortedCharacter_10,
  output [8:0]  io_outputs_sortedCharacter_11,
  output [8:0]  io_outputs_sortedCharacter_12,
  output [8:0]  io_outputs_sortedCharacter_13,
  output [8:0]  io_outputs_sortedCharacter_14,
  output [8:0]  io_outputs_sortedCharacter_15,
  output [8:0]  io_outputs_sortedCharacter_16,
  output [8:0]  io_outputs_sortedCharacter_17,
  output [8:0]  io_outputs_sortedCharacter_18,
  output [8:0]  io_outputs_sortedCharacter_19,
  output [8:0]  io_outputs_sortedCharacter_20,
  output [8:0]  io_outputs_sortedCharacter_21,
  output [8:0]  io_outputs_sortedCharacter_22,
  output [8:0]  io_outputs_sortedCharacter_23,
  output [8:0]  io_outputs_sortedCharacter_24,
  output [8:0]  io_outputs_sortedCharacter_25,
  output [8:0]  io_outputs_sortedCharacter_26,
  output [8:0]  io_outputs_sortedCharacter_27,
  output [8:0]  io_outputs_sortedCharacter_28,
  output [8:0]  io_outputs_sortedCharacter_29,
  output [8:0]  io_outputs_sortedCharacter_30,
  output [8:0]  io_outputs_sortedCharacter_31,
  output        io_finished
);
  wire [11:0] input__io_input_currentByteOut; // @[characterFrequencyModule.scala 24:21]
  wire [7:0] input__io_input_dataIn_0; // @[characterFrequencyModule.scala 24:21]
  wire  input__io_input_valid; // @[characterFrequencyModule.scala 24:21]
  wire  input__io_input_ready; // @[characterFrequencyModule.scala 24:21]
  wire [11:0] input__io_currentByte; // @[characterFrequencyModule.scala 24:21]
  wire  input__io_dataOut_ready; // @[characterFrequencyModule.scala 24:21]
  wire  input__io_dataOut_valid; // @[characterFrequencyModule.scala 24:21]
  wire [7:0] input__io_dataOut_bits_0; // @[characterFrequencyModule.scala 24:21]
  wire  count_clock; // @[characterFrequencyModule.scala 26:21]
  wire  count_reset; // @[characterFrequencyModule.scala 26:21]
  wire  count_io_start; // @[characterFrequencyModule.scala 26:21]
  wire  count_io_dataIn_ready; // @[characterFrequencyModule.scala 26:21]
  wire [7:0] count_io_dataIn_bits_0; // @[characterFrequencyModule.scala 26:21]
  wire [11:0] count_io_currentByte; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_0; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_1; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_2; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_3; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_4; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_5; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_6; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_7; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_8; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_9; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_10; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_11; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_12; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_13; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_14; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_15; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_16; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_17; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_18; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_19; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_20; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_21; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_22; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_23; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_24; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_25; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_26; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_27; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_28; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_29; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_30; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_31; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_32; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_33; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_34; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_35; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_36; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_37; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_38; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_39; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_40; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_41; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_42; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_43; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_44; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_45; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_46; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_47; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_48; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_49; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_50; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_51; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_52; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_53; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_54; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_55; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_56; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_57; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_58; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_59; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_60; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_61; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_62; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_63; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_64; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_65; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_66; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_67; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_68; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_69; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_70; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_71; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_72; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_73; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_74; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_75; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_76; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_77; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_78; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_79; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_80; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_81; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_82; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_83; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_84; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_85; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_86; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_87; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_88; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_89; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_90; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_91; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_92; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_93; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_94; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_95; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_96; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_97; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_98; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_99; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_100; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_101; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_102; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_103; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_104; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_105; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_106; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_107; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_108; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_109; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_110; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_111; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_112; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_113; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_114; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_115; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_116; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_117; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_118; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_119; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_120; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_121; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_122; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_123; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_124; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_125; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_126; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_127; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_128; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_129; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_130; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_131; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_132; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_133; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_134; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_135; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_136; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_137; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_138; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_139; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_140; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_141; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_142; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_143; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_144; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_145; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_146; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_147; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_148; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_149; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_150; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_151; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_152; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_153; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_154; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_155; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_156; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_157; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_158; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_159; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_160; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_161; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_162; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_163; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_164; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_165; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_166; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_167; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_168; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_169; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_170; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_171; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_172; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_173; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_174; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_175; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_176; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_177; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_178; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_179; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_180; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_181; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_182; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_183; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_184; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_185; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_186; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_187; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_188; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_189; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_190; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_191; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_192; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_193; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_194; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_195; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_196; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_197; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_198; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_199; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_200; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_201; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_202; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_203; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_204; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_205; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_206; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_207; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_208; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_209; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_210; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_211; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_212; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_213; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_214; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_215; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_216; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_217; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_218; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_219; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_220; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_221; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_222; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_223; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_224; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_225; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_226; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_227; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_228; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_229; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_230; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_231; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_232; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_233; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_234; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_235; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_236; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_237; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_238; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_239; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_240; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_241; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_242; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_243; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_244; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_245; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_246; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_247; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_248; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_249; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_250; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_251; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_252; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_253; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_254; // @[characterFrequencyModule.scala 26:21]
  wire [12:0] count_io_frequencies_255; // @[characterFrequencyModule.scala 26:21]
  wire  count_io_finished; // @[characterFrequencyModule.scala 26:21]
  wire  sort_clock; // @[characterFrequencyModule.scala 28:20]
  wire  sort_reset; // @[characterFrequencyModule.scala 28:20]
  wire  sort_io_start; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_0; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_1; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_2; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_3; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_4; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_5; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_6; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_7; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_8; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_9; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_10; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_11; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_12; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_13; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_14; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_15; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_16; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_17; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_18; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_19; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_20; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_21; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_22; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_23; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_24; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_25; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_26; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_27; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_28; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_29; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_30; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_31; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_32; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_33; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_34; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_35; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_36; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_37; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_38; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_39; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_40; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_41; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_42; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_43; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_44; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_45; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_46; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_47; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_48; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_49; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_50; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_51; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_52; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_53; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_54; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_55; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_56; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_57; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_58; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_59; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_60; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_61; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_62; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_63; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_64; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_65; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_66; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_67; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_68; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_69; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_70; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_71; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_72; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_73; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_74; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_75; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_76; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_77; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_78; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_79; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_80; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_81; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_82; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_83; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_84; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_85; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_86; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_87; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_88; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_89; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_90; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_91; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_92; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_93; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_94; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_95; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_96; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_97; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_98; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_99; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_100; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_101; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_102; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_103; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_104; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_105; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_106; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_107; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_108; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_109; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_110; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_111; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_112; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_113; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_114; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_115; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_116; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_117; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_118; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_119; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_120; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_121; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_122; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_123; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_124; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_125; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_126; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_127; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_128; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_129; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_130; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_131; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_132; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_133; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_134; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_135; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_136; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_137; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_138; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_139; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_140; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_141; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_142; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_143; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_144; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_145; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_146; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_147; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_148; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_149; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_150; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_151; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_152; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_153; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_154; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_155; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_156; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_157; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_158; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_159; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_160; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_161; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_162; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_163; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_164; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_165; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_166; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_167; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_168; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_169; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_170; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_171; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_172; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_173; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_174; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_175; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_176; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_177; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_178; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_179; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_180; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_181; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_182; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_183; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_184; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_185; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_186; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_187; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_188; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_189; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_190; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_191; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_192; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_193; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_194; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_195; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_196; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_197; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_198; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_199; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_200; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_201; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_202; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_203; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_204; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_205; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_206; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_207; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_208; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_209; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_210; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_211; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_212; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_213; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_214; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_215; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_216; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_217; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_218; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_219; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_220; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_221; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_222; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_223; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_224; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_225; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_226; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_227; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_228; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_229; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_230; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_231; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_232; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_233; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_234; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_235; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_236; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_237; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_238; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_239; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_240; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_241; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_242; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_243; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_244; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_245; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_246; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_247; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_248; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_249; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_250; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_251; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_252; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_253; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_254; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_dataIn_255; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_0; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_1; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_2; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_3; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_4; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_5; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_6; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_7; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_8; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_9; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_10; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_11; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_12; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_13; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_14; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_15; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_16; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_17; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_18; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_19; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_20; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_21; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_22; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_23; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_24; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_25; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_26; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_27; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_28; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_29; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_30; // @[characterFrequencyModule.scala 28:20]
  wire [12:0] sort_io_sortedFrequency_31; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_0; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_1; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_2; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_3; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_4; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_5; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_6; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_7; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_8; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_9; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_10; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_11; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_12; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_13; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_14; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_15; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_16; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_17; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_18; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_19; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_20; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_21; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_22; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_23; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_24; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_25; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_26; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_27; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_28; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_29; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_30; // @[characterFrequencyModule.scala 28:20]
  wire [8:0] sort_io_sortedCharacter_31; // @[characterFrequencyModule.scala 28:20]
  wire  sort_io_finished; // @[characterFrequencyModule.scala 28:20]
  reg  previousCountFinished; // @[characterFrequencyModule.scala 32:38]
  reg [31:0] _RAND_0;
  wire  _T = ~previousCountFinished; // @[characterFrequencyModule.scala 38:41]
  compressorInput input_ ( // @[characterFrequencyModule.scala 24:21]
    .io_input_currentByteOut(input__io_input_currentByteOut),
    .io_input_dataIn_0(input__io_input_dataIn_0),
    .io_input_valid(input__io_input_valid),
    .io_input_ready(input__io_input_ready),
    .io_currentByte(input__io_currentByte),
    .io_dataOut_ready(input__io_dataOut_ready),
    .io_dataOut_valid(input__io_dataOut_valid),
    .io_dataOut_bits_0(input__io_dataOut_bits_0)
  );
  characterFrequencyCounter count ( // @[characterFrequencyModule.scala 26:21]
    .clock(count_clock),
    .reset(count_reset),
    .io_start(count_io_start),
    .io_dataIn_ready(count_io_dataIn_ready),
    .io_dataIn_bits_0(count_io_dataIn_bits_0),
    .io_currentByte(count_io_currentByte),
    .io_frequencies_0(count_io_frequencies_0),
    .io_frequencies_1(count_io_frequencies_1),
    .io_frequencies_2(count_io_frequencies_2),
    .io_frequencies_3(count_io_frequencies_3),
    .io_frequencies_4(count_io_frequencies_4),
    .io_frequencies_5(count_io_frequencies_5),
    .io_frequencies_6(count_io_frequencies_6),
    .io_frequencies_7(count_io_frequencies_7),
    .io_frequencies_8(count_io_frequencies_8),
    .io_frequencies_9(count_io_frequencies_9),
    .io_frequencies_10(count_io_frequencies_10),
    .io_frequencies_11(count_io_frequencies_11),
    .io_frequencies_12(count_io_frequencies_12),
    .io_frequencies_13(count_io_frequencies_13),
    .io_frequencies_14(count_io_frequencies_14),
    .io_frequencies_15(count_io_frequencies_15),
    .io_frequencies_16(count_io_frequencies_16),
    .io_frequencies_17(count_io_frequencies_17),
    .io_frequencies_18(count_io_frequencies_18),
    .io_frequencies_19(count_io_frequencies_19),
    .io_frequencies_20(count_io_frequencies_20),
    .io_frequencies_21(count_io_frequencies_21),
    .io_frequencies_22(count_io_frequencies_22),
    .io_frequencies_23(count_io_frequencies_23),
    .io_frequencies_24(count_io_frequencies_24),
    .io_frequencies_25(count_io_frequencies_25),
    .io_frequencies_26(count_io_frequencies_26),
    .io_frequencies_27(count_io_frequencies_27),
    .io_frequencies_28(count_io_frequencies_28),
    .io_frequencies_29(count_io_frequencies_29),
    .io_frequencies_30(count_io_frequencies_30),
    .io_frequencies_31(count_io_frequencies_31),
    .io_frequencies_32(count_io_frequencies_32),
    .io_frequencies_33(count_io_frequencies_33),
    .io_frequencies_34(count_io_frequencies_34),
    .io_frequencies_35(count_io_frequencies_35),
    .io_frequencies_36(count_io_frequencies_36),
    .io_frequencies_37(count_io_frequencies_37),
    .io_frequencies_38(count_io_frequencies_38),
    .io_frequencies_39(count_io_frequencies_39),
    .io_frequencies_40(count_io_frequencies_40),
    .io_frequencies_41(count_io_frequencies_41),
    .io_frequencies_42(count_io_frequencies_42),
    .io_frequencies_43(count_io_frequencies_43),
    .io_frequencies_44(count_io_frequencies_44),
    .io_frequencies_45(count_io_frequencies_45),
    .io_frequencies_46(count_io_frequencies_46),
    .io_frequencies_47(count_io_frequencies_47),
    .io_frequencies_48(count_io_frequencies_48),
    .io_frequencies_49(count_io_frequencies_49),
    .io_frequencies_50(count_io_frequencies_50),
    .io_frequencies_51(count_io_frequencies_51),
    .io_frequencies_52(count_io_frequencies_52),
    .io_frequencies_53(count_io_frequencies_53),
    .io_frequencies_54(count_io_frequencies_54),
    .io_frequencies_55(count_io_frequencies_55),
    .io_frequencies_56(count_io_frequencies_56),
    .io_frequencies_57(count_io_frequencies_57),
    .io_frequencies_58(count_io_frequencies_58),
    .io_frequencies_59(count_io_frequencies_59),
    .io_frequencies_60(count_io_frequencies_60),
    .io_frequencies_61(count_io_frequencies_61),
    .io_frequencies_62(count_io_frequencies_62),
    .io_frequencies_63(count_io_frequencies_63),
    .io_frequencies_64(count_io_frequencies_64),
    .io_frequencies_65(count_io_frequencies_65),
    .io_frequencies_66(count_io_frequencies_66),
    .io_frequencies_67(count_io_frequencies_67),
    .io_frequencies_68(count_io_frequencies_68),
    .io_frequencies_69(count_io_frequencies_69),
    .io_frequencies_70(count_io_frequencies_70),
    .io_frequencies_71(count_io_frequencies_71),
    .io_frequencies_72(count_io_frequencies_72),
    .io_frequencies_73(count_io_frequencies_73),
    .io_frequencies_74(count_io_frequencies_74),
    .io_frequencies_75(count_io_frequencies_75),
    .io_frequencies_76(count_io_frequencies_76),
    .io_frequencies_77(count_io_frequencies_77),
    .io_frequencies_78(count_io_frequencies_78),
    .io_frequencies_79(count_io_frequencies_79),
    .io_frequencies_80(count_io_frequencies_80),
    .io_frequencies_81(count_io_frequencies_81),
    .io_frequencies_82(count_io_frequencies_82),
    .io_frequencies_83(count_io_frequencies_83),
    .io_frequencies_84(count_io_frequencies_84),
    .io_frequencies_85(count_io_frequencies_85),
    .io_frequencies_86(count_io_frequencies_86),
    .io_frequencies_87(count_io_frequencies_87),
    .io_frequencies_88(count_io_frequencies_88),
    .io_frequencies_89(count_io_frequencies_89),
    .io_frequencies_90(count_io_frequencies_90),
    .io_frequencies_91(count_io_frequencies_91),
    .io_frequencies_92(count_io_frequencies_92),
    .io_frequencies_93(count_io_frequencies_93),
    .io_frequencies_94(count_io_frequencies_94),
    .io_frequencies_95(count_io_frequencies_95),
    .io_frequencies_96(count_io_frequencies_96),
    .io_frequencies_97(count_io_frequencies_97),
    .io_frequencies_98(count_io_frequencies_98),
    .io_frequencies_99(count_io_frequencies_99),
    .io_frequencies_100(count_io_frequencies_100),
    .io_frequencies_101(count_io_frequencies_101),
    .io_frequencies_102(count_io_frequencies_102),
    .io_frequencies_103(count_io_frequencies_103),
    .io_frequencies_104(count_io_frequencies_104),
    .io_frequencies_105(count_io_frequencies_105),
    .io_frequencies_106(count_io_frequencies_106),
    .io_frequencies_107(count_io_frequencies_107),
    .io_frequencies_108(count_io_frequencies_108),
    .io_frequencies_109(count_io_frequencies_109),
    .io_frequencies_110(count_io_frequencies_110),
    .io_frequencies_111(count_io_frequencies_111),
    .io_frequencies_112(count_io_frequencies_112),
    .io_frequencies_113(count_io_frequencies_113),
    .io_frequencies_114(count_io_frequencies_114),
    .io_frequencies_115(count_io_frequencies_115),
    .io_frequencies_116(count_io_frequencies_116),
    .io_frequencies_117(count_io_frequencies_117),
    .io_frequencies_118(count_io_frequencies_118),
    .io_frequencies_119(count_io_frequencies_119),
    .io_frequencies_120(count_io_frequencies_120),
    .io_frequencies_121(count_io_frequencies_121),
    .io_frequencies_122(count_io_frequencies_122),
    .io_frequencies_123(count_io_frequencies_123),
    .io_frequencies_124(count_io_frequencies_124),
    .io_frequencies_125(count_io_frequencies_125),
    .io_frequencies_126(count_io_frequencies_126),
    .io_frequencies_127(count_io_frequencies_127),
    .io_frequencies_128(count_io_frequencies_128),
    .io_frequencies_129(count_io_frequencies_129),
    .io_frequencies_130(count_io_frequencies_130),
    .io_frequencies_131(count_io_frequencies_131),
    .io_frequencies_132(count_io_frequencies_132),
    .io_frequencies_133(count_io_frequencies_133),
    .io_frequencies_134(count_io_frequencies_134),
    .io_frequencies_135(count_io_frequencies_135),
    .io_frequencies_136(count_io_frequencies_136),
    .io_frequencies_137(count_io_frequencies_137),
    .io_frequencies_138(count_io_frequencies_138),
    .io_frequencies_139(count_io_frequencies_139),
    .io_frequencies_140(count_io_frequencies_140),
    .io_frequencies_141(count_io_frequencies_141),
    .io_frequencies_142(count_io_frequencies_142),
    .io_frequencies_143(count_io_frequencies_143),
    .io_frequencies_144(count_io_frequencies_144),
    .io_frequencies_145(count_io_frequencies_145),
    .io_frequencies_146(count_io_frequencies_146),
    .io_frequencies_147(count_io_frequencies_147),
    .io_frequencies_148(count_io_frequencies_148),
    .io_frequencies_149(count_io_frequencies_149),
    .io_frequencies_150(count_io_frequencies_150),
    .io_frequencies_151(count_io_frequencies_151),
    .io_frequencies_152(count_io_frequencies_152),
    .io_frequencies_153(count_io_frequencies_153),
    .io_frequencies_154(count_io_frequencies_154),
    .io_frequencies_155(count_io_frequencies_155),
    .io_frequencies_156(count_io_frequencies_156),
    .io_frequencies_157(count_io_frequencies_157),
    .io_frequencies_158(count_io_frequencies_158),
    .io_frequencies_159(count_io_frequencies_159),
    .io_frequencies_160(count_io_frequencies_160),
    .io_frequencies_161(count_io_frequencies_161),
    .io_frequencies_162(count_io_frequencies_162),
    .io_frequencies_163(count_io_frequencies_163),
    .io_frequencies_164(count_io_frequencies_164),
    .io_frequencies_165(count_io_frequencies_165),
    .io_frequencies_166(count_io_frequencies_166),
    .io_frequencies_167(count_io_frequencies_167),
    .io_frequencies_168(count_io_frequencies_168),
    .io_frequencies_169(count_io_frequencies_169),
    .io_frequencies_170(count_io_frequencies_170),
    .io_frequencies_171(count_io_frequencies_171),
    .io_frequencies_172(count_io_frequencies_172),
    .io_frequencies_173(count_io_frequencies_173),
    .io_frequencies_174(count_io_frequencies_174),
    .io_frequencies_175(count_io_frequencies_175),
    .io_frequencies_176(count_io_frequencies_176),
    .io_frequencies_177(count_io_frequencies_177),
    .io_frequencies_178(count_io_frequencies_178),
    .io_frequencies_179(count_io_frequencies_179),
    .io_frequencies_180(count_io_frequencies_180),
    .io_frequencies_181(count_io_frequencies_181),
    .io_frequencies_182(count_io_frequencies_182),
    .io_frequencies_183(count_io_frequencies_183),
    .io_frequencies_184(count_io_frequencies_184),
    .io_frequencies_185(count_io_frequencies_185),
    .io_frequencies_186(count_io_frequencies_186),
    .io_frequencies_187(count_io_frequencies_187),
    .io_frequencies_188(count_io_frequencies_188),
    .io_frequencies_189(count_io_frequencies_189),
    .io_frequencies_190(count_io_frequencies_190),
    .io_frequencies_191(count_io_frequencies_191),
    .io_frequencies_192(count_io_frequencies_192),
    .io_frequencies_193(count_io_frequencies_193),
    .io_frequencies_194(count_io_frequencies_194),
    .io_frequencies_195(count_io_frequencies_195),
    .io_frequencies_196(count_io_frequencies_196),
    .io_frequencies_197(count_io_frequencies_197),
    .io_frequencies_198(count_io_frequencies_198),
    .io_frequencies_199(count_io_frequencies_199),
    .io_frequencies_200(count_io_frequencies_200),
    .io_frequencies_201(count_io_frequencies_201),
    .io_frequencies_202(count_io_frequencies_202),
    .io_frequencies_203(count_io_frequencies_203),
    .io_frequencies_204(count_io_frequencies_204),
    .io_frequencies_205(count_io_frequencies_205),
    .io_frequencies_206(count_io_frequencies_206),
    .io_frequencies_207(count_io_frequencies_207),
    .io_frequencies_208(count_io_frequencies_208),
    .io_frequencies_209(count_io_frequencies_209),
    .io_frequencies_210(count_io_frequencies_210),
    .io_frequencies_211(count_io_frequencies_211),
    .io_frequencies_212(count_io_frequencies_212),
    .io_frequencies_213(count_io_frequencies_213),
    .io_frequencies_214(count_io_frequencies_214),
    .io_frequencies_215(count_io_frequencies_215),
    .io_frequencies_216(count_io_frequencies_216),
    .io_frequencies_217(count_io_frequencies_217),
    .io_frequencies_218(count_io_frequencies_218),
    .io_frequencies_219(count_io_frequencies_219),
    .io_frequencies_220(count_io_frequencies_220),
    .io_frequencies_221(count_io_frequencies_221),
    .io_frequencies_222(count_io_frequencies_222),
    .io_frequencies_223(count_io_frequencies_223),
    .io_frequencies_224(count_io_frequencies_224),
    .io_frequencies_225(count_io_frequencies_225),
    .io_frequencies_226(count_io_frequencies_226),
    .io_frequencies_227(count_io_frequencies_227),
    .io_frequencies_228(count_io_frequencies_228),
    .io_frequencies_229(count_io_frequencies_229),
    .io_frequencies_230(count_io_frequencies_230),
    .io_frequencies_231(count_io_frequencies_231),
    .io_frequencies_232(count_io_frequencies_232),
    .io_frequencies_233(count_io_frequencies_233),
    .io_frequencies_234(count_io_frequencies_234),
    .io_frequencies_235(count_io_frequencies_235),
    .io_frequencies_236(count_io_frequencies_236),
    .io_frequencies_237(count_io_frequencies_237),
    .io_frequencies_238(count_io_frequencies_238),
    .io_frequencies_239(count_io_frequencies_239),
    .io_frequencies_240(count_io_frequencies_240),
    .io_frequencies_241(count_io_frequencies_241),
    .io_frequencies_242(count_io_frequencies_242),
    .io_frequencies_243(count_io_frequencies_243),
    .io_frequencies_244(count_io_frequencies_244),
    .io_frequencies_245(count_io_frequencies_245),
    .io_frequencies_246(count_io_frequencies_246),
    .io_frequencies_247(count_io_frequencies_247),
    .io_frequencies_248(count_io_frequencies_248),
    .io_frequencies_249(count_io_frequencies_249),
    .io_frequencies_250(count_io_frequencies_250),
    .io_frequencies_251(count_io_frequencies_251),
    .io_frequencies_252(count_io_frequencies_252),
    .io_frequencies_253(count_io_frequencies_253),
    .io_frequencies_254(count_io_frequencies_254),
    .io_frequencies_255(count_io_frequencies_255),
    .io_finished(count_io_finished)
  );
  characterFrequencySort sort ( // @[characterFrequencyModule.scala 28:20]
    .clock(sort_clock),
    .reset(sort_reset),
    .io_start(sort_io_start),
    .io_dataIn_0(sort_io_dataIn_0),
    .io_dataIn_1(sort_io_dataIn_1),
    .io_dataIn_2(sort_io_dataIn_2),
    .io_dataIn_3(sort_io_dataIn_3),
    .io_dataIn_4(sort_io_dataIn_4),
    .io_dataIn_5(sort_io_dataIn_5),
    .io_dataIn_6(sort_io_dataIn_6),
    .io_dataIn_7(sort_io_dataIn_7),
    .io_dataIn_8(sort_io_dataIn_8),
    .io_dataIn_9(sort_io_dataIn_9),
    .io_dataIn_10(sort_io_dataIn_10),
    .io_dataIn_11(sort_io_dataIn_11),
    .io_dataIn_12(sort_io_dataIn_12),
    .io_dataIn_13(sort_io_dataIn_13),
    .io_dataIn_14(sort_io_dataIn_14),
    .io_dataIn_15(sort_io_dataIn_15),
    .io_dataIn_16(sort_io_dataIn_16),
    .io_dataIn_17(sort_io_dataIn_17),
    .io_dataIn_18(sort_io_dataIn_18),
    .io_dataIn_19(sort_io_dataIn_19),
    .io_dataIn_20(sort_io_dataIn_20),
    .io_dataIn_21(sort_io_dataIn_21),
    .io_dataIn_22(sort_io_dataIn_22),
    .io_dataIn_23(sort_io_dataIn_23),
    .io_dataIn_24(sort_io_dataIn_24),
    .io_dataIn_25(sort_io_dataIn_25),
    .io_dataIn_26(sort_io_dataIn_26),
    .io_dataIn_27(sort_io_dataIn_27),
    .io_dataIn_28(sort_io_dataIn_28),
    .io_dataIn_29(sort_io_dataIn_29),
    .io_dataIn_30(sort_io_dataIn_30),
    .io_dataIn_31(sort_io_dataIn_31),
    .io_dataIn_32(sort_io_dataIn_32),
    .io_dataIn_33(sort_io_dataIn_33),
    .io_dataIn_34(sort_io_dataIn_34),
    .io_dataIn_35(sort_io_dataIn_35),
    .io_dataIn_36(sort_io_dataIn_36),
    .io_dataIn_37(sort_io_dataIn_37),
    .io_dataIn_38(sort_io_dataIn_38),
    .io_dataIn_39(sort_io_dataIn_39),
    .io_dataIn_40(sort_io_dataIn_40),
    .io_dataIn_41(sort_io_dataIn_41),
    .io_dataIn_42(sort_io_dataIn_42),
    .io_dataIn_43(sort_io_dataIn_43),
    .io_dataIn_44(sort_io_dataIn_44),
    .io_dataIn_45(sort_io_dataIn_45),
    .io_dataIn_46(sort_io_dataIn_46),
    .io_dataIn_47(sort_io_dataIn_47),
    .io_dataIn_48(sort_io_dataIn_48),
    .io_dataIn_49(sort_io_dataIn_49),
    .io_dataIn_50(sort_io_dataIn_50),
    .io_dataIn_51(sort_io_dataIn_51),
    .io_dataIn_52(sort_io_dataIn_52),
    .io_dataIn_53(sort_io_dataIn_53),
    .io_dataIn_54(sort_io_dataIn_54),
    .io_dataIn_55(sort_io_dataIn_55),
    .io_dataIn_56(sort_io_dataIn_56),
    .io_dataIn_57(sort_io_dataIn_57),
    .io_dataIn_58(sort_io_dataIn_58),
    .io_dataIn_59(sort_io_dataIn_59),
    .io_dataIn_60(sort_io_dataIn_60),
    .io_dataIn_61(sort_io_dataIn_61),
    .io_dataIn_62(sort_io_dataIn_62),
    .io_dataIn_63(sort_io_dataIn_63),
    .io_dataIn_64(sort_io_dataIn_64),
    .io_dataIn_65(sort_io_dataIn_65),
    .io_dataIn_66(sort_io_dataIn_66),
    .io_dataIn_67(sort_io_dataIn_67),
    .io_dataIn_68(sort_io_dataIn_68),
    .io_dataIn_69(sort_io_dataIn_69),
    .io_dataIn_70(sort_io_dataIn_70),
    .io_dataIn_71(sort_io_dataIn_71),
    .io_dataIn_72(sort_io_dataIn_72),
    .io_dataIn_73(sort_io_dataIn_73),
    .io_dataIn_74(sort_io_dataIn_74),
    .io_dataIn_75(sort_io_dataIn_75),
    .io_dataIn_76(sort_io_dataIn_76),
    .io_dataIn_77(sort_io_dataIn_77),
    .io_dataIn_78(sort_io_dataIn_78),
    .io_dataIn_79(sort_io_dataIn_79),
    .io_dataIn_80(sort_io_dataIn_80),
    .io_dataIn_81(sort_io_dataIn_81),
    .io_dataIn_82(sort_io_dataIn_82),
    .io_dataIn_83(sort_io_dataIn_83),
    .io_dataIn_84(sort_io_dataIn_84),
    .io_dataIn_85(sort_io_dataIn_85),
    .io_dataIn_86(sort_io_dataIn_86),
    .io_dataIn_87(sort_io_dataIn_87),
    .io_dataIn_88(sort_io_dataIn_88),
    .io_dataIn_89(sort_io_dataIn_89),
    .io_dataIn_90(sort_io_dataIn_90),
    .io_dataIn_91(sort_io_dataIn_91),
    .io_dataIn_92(sort_io_dataIn_92),
    .io_dataIn_93(sort_io_dataIn_93),
    .io_dataIn_94(sort_io_dataIn_94),
    .io_dataIn_95(sort_io_dataIn_95),
    .io_dataIn_96(sort_io_dataIn_96),
    .io_dataIn_97(sort_io_dataIn_97),
    .io_dataIn_98(sort_io_dataIn_98),
    .io_dataIn_99(sort_io_dataIn_99),
    .io_dataIn_100(sort_io_dataIn_100),
    .io_dataIn_101(sort_io_dataIn_101),
    .io_dataIn_102(sort_io_dataIn_102),
    .io_dataIn_103(sort_io_dataIn_103),
    .io_dataIn_104(sort_io_dataIn_104),
    .io_dataIn_105(sort_io_dataIn_105),
    .io_dataIn_106(sort_io_dataIn_106),
    .io_dataIn_107(sort_io_dataIn_107),
    .io_dataIn_108(sort_io_dataIn_108),
    .io_dataIn_109(sort_io_dataIn_109),
    .io_dataIn_110(sort_io_dataIn_110),
    .io_dataIn_111(sort_io_dataIn_111),
    .io_dataIn_112(sort_io_dataIn_112),
    .io_dataIn_113(sort_io_dataIn_113),
    .io_dataIn_114(sort_io_dataIn_114),
    .io_dataIn_115(sort_io_dataIn_115),
    .io_dataIn_116(sort_io_dataIn_116),
    .io_dataIn_117(sort_io_dataIn_117),
    .io_dataIn_118(sort_io_dataIn_118),
    .io_dataIn_119(sort_io_dataIn_119),
    .io_dataIn_120(sort_io_dataIn_120),
    .io_dataIn_121(sort_io_dataIn_121),
    .io_dataIn_122(sort_io_dataIn_122),
    .io_dataIn_123(sort_io_dataIn_123),
    .io_dataIn_124(sort_io_dataIn_124),
    .io_dataIn_125(sort_io_dataIn_125),
    .io_dataIn_126(sort_io_dataIn_126),
    .io_dataIn_127(sort_io_dataIn_127),
    .io_dataIn_128(sort_io_dataIn_128),
    .io_dataIn_129(sort_io_dataIn_129),
    .io_dataIn_130(sort_io_dataIn_130),
    .io_dataIn_131(sort_io_dataIn_131),
    .io_dataIn_132(sort_io_dataIn_132),
    .io_dataIn_133(sort_io_dataIn_133),
    .io_dataIn_134(sort_io_dataIn_134),
    .io_dataIn_135(sort_io_dataIn_135),
    .io_dataIn_136(sort_io_dataIn_136),
    .io_dataIn_137(sort_io_dataIn_137),
    .io_dataIn_138(sort_io_dataIn_138),
    .io_dataIn_139(sort_io_dataIn_139),
    .io_dataIn_140(sort_io_dataIn_140),
    .io_dataIn_141(sort_io_dataIn_141),
    .io_dataIn_142(sort_io_dataIn_142),
    .io_dataIn_143(sort_io_dataIn_143),
    .io_dataIn_144(sort_io_dataIn_144),
    .io_dataIn_145(sort_io_dataIn_145),
    .io_dataIn_146(sort_io_dataIn_146),
    .io_dataIn_147(sort_io_dataIn_147),
    .io_dataIn_148(sort_io_dataIn_148),
    .io_dataIn_149(sort_io_dataIn_149),
    .io_dataIn_150(sort_io_dataIn_150),
    .io_dataIn_151(sort_io_dataIn_151),
    .io_dataIn_152(sort_io_dataIn_152),
    .io_dataIn_153(sort_io_dataIn_153),
    .io_dataIn_154(sort_io_dataIn_154),
    .io_dataIn_155(sort_io_dataIn_155),
    .io_dataIn_156(sort_io_dataIn_156),
    .io_dataIn_157(sort_io_dataIn_157),
    .io_dataIn_158(sort_io_dataIn_158),
    .io_dataIn_159(sort_io_dataIn_159),
    .io_dataIn_160(sort_io_dataIn_160),
    .io_dataIn_161(sort_io_dataIn_161),
    .io_dataIn_162(sort_io_dataIn_162),
    .io_dataIn_163(sort_io_dataIn_163),
    .io_dataIn_164(sort_io_dataIn_164),
    .io_dataIn_165(sort_io_dataIn_165),
    .io_dataIn_166(sort_io_dataIn_166),
    .io_dataIn_167(sort_io_dataIn_167),
    .io_dataIn_168(sort_io_dataIn_168),
    .io_dataIn_169(sort_io_dataIn_169),
    .io_dataIn_170(sort_io_dataIn_170),
    .io_dataIn_171(sort_io_dataIn_171),
    .io_dataIn_172(sort_io_dataIn_172),
    .io_dataIn_173(sort_io_dataIn_173),
    .io_dataIn_174(sort_io_dataIn_174),
    .io_dataIn_175(sort_io_dataIn_175),
    .io_dataIn_176(sort_io_dataIn_176),
    .io_dataIn_177(sort_io_dataIn_177),
    .io_dataIn_178(sort_io_dataIn_178),
    .io_dataIn_179(sort_io_dataIn_179),
    .io_dataIn_180(sort_io_dataIn_180),
    .io_dataIn_181(sort_io_dataIn_181),
    .io_dataIn_182(sort_io_dataIn_182),
    .io_dataIn_183(sort_io_dataIn_183),
    .io_dataIn_184(sort_io_dataIn_184),
    .io_dataIn_185(sort_io_dataIn_185),
    .io_dataIn_186(sort_io_dataIn_186),
    .io_dataIn_187(sort_io_dataIn_187),
    .io_dataIn_188(sort_io_dataIn_188),
    .io_dataIn_189(sort_io_dataIn_189),
    .io_dataIn_190(sort_io_dataIn_190),
    .io_dataIn_191(sort_io_dataIn_191),
    .io_dataIn_192(sort_io_dataIn_192),
    .io_dataIn_193(sort_io_dataIn_193),
    .io_dataIn_194(sort_io_dataIn_194),
    .io_dataIn_195(sort_io_dataIn_195),
    .io_dataIn_196(sort_io_dataIn_196),
    .io_dataIn_197(sort_io_dataIn_197),
    .io_dataIn_198(sort_io_dataIn_198),
    .io_dataIn_199(sort_io_dataIn_199),
    .io_dataIn_200(sort_io_dataIn_200),
    .io_dataIn_201(sort_io_dataIn_201),
    .io_dataIn_202(sort_io_dataIn_202),
    .io_dataIn_203(sort_io_dataIn_203),
    .io_dataIn_204(sort_io_dataIn_204),
    .io_dataIn_205(sort_io_dataIn_205),
    .io_dataIn_206(sort_io_dataIn_206),
    .io_dataIn_207(sort_io_dataIn_207),
    .io_dataIn_208(sort_io_dataIn_208),
    .io_dataIn_209(sort_io_dataIn_209),
    .io_dataIn_210(sort_io_dataIn_210),
    .io_dataIn_211(sort_io_dataIn_211),
    .io_dataIn_212(sort_io_dataIn_212),
    .io_dataIn_213(sort_io_dataIn_213),
    .io_dataIn_214(sort_io_dataIn_214),
    .io_dataIn_215(sort_io_dataIn_215),
    .io_dataIn_216(sort_io_dataIn_216),
    .io_dataIn_217(sort_io_dataIn_217),
    .io_dataIn_218(sort_io_dataIn_218),
    .io_dataIn_219(sort_io_dataIn_219),
    .io_dataIn_220(sort_io_dataIn_220),
    .io_dataIn_221(sort_io_dataIn_221),
    .io_dataIn_222(sort_io_dataIn_222),
    .io_dataIn_223(sort_io_dataIn_223),
    .io_dataIn_224(sort_io_dataIn_224),
    .io_dataIn_225(sort_io_dataIn_225),
    .io_dataIn_226(sort_io_dataIn_226),
    .io_dataIn_227(sort_io_dataIn_227),
    .io_dataIn_228(sort_io_dataIn_228),
    .io_dataIn_229(sort_io_dataIn_229),
    .io_dataIn_230(sort_io_dataIn_230),
    .io_dataIn_231(sort_io_dataIn_231),
    .io_dataIn_232(sort_io_dataIn_232),
    .io_dataIn_233(sort_io_dataIn_233),
    .io_dataIn_234(sort_io_dataIn_234),
    .io_dataIn_235(sort_io_dataIn_235),
    .io_dataIn_236(sort_io_dataIn_236),
    .io_dataIn_237(sort_io_dataIn_237),
    .io_dataIn_238(sort_io_dataIn_238),
    .io_dataIn_239(sort_io_dataIn_239),
    .io_dataIn_240(sort_io_dataIn_240),
    .io_dataIn_241(sort_io_dataIn_241),
    .io_dataIn_242(sort_io_dataIn_242),
    .io_dataIn_243(sort_io_dataIn_243),
    .io_dataIn_244(sort_io_dataIn_244),
    .io_dataIn_245(sort_io_dataIn_245),
    .io_dataIn_246(sort_io_dataIn_246),
    .io_dataIn_247(sort_io_dataIn_247),
    .io_dataIn_248(sort_io_dataIn_248),
    .io_dataIn_249(sort_io_dataIn_249),
    .io_dataIn_250(sort_io_dataIn_250),
    .io_dataIn_251(sort_io_dataIn_251),
    .io_dataIn_252(sort_io_dataIn_252),
    .io_dataIn_253(sort_io_dataIn_253),
    .io_dataIn_254(sort_io_dataIn_254),
    .io_dataIn_255(sort_io_dataIn_255),
    .io_sortedFrequency_0(sort_io_sortedFrequency_0),
    .io_sortedFrequency_1(sort_io_sortedFrequency_1),
    .io_sortedFrequency_2(sort_io_sortedFrequency_2),
    .io_sortedFrequency_3(sort_io_sortedFrequency_3),
    .io_sortedFrequency_4(sort_io_sortedFrequency_4),
    .io_sortedFrequency_5(sort_io_sortedFrequency_5),
    .io_sortedFrequency_6(sort_io_sortedFrequency_6),
    .io_sortedFrequency_7(sort_io_sortedFrequency_7),
    .io_sortedFrequency_8(sort_io_sortedFrequency_8),
    .io_sortedFrequency_9(sort_io_sortedFrequency_9),
    .io_sortedFrequency_10(sort_io_sortedFrequency_10),
    .io_sortedFrequency_11(sort_io_sortedFrequency_11),
    .io_sortedFrequency_12(sort_io_sortedFrequency_12),
    .io_sortedFrequency_13(sort_io_sortedFrequency_13),
    .io_sortedFrequency_14(sort_io_sortedFrequency_14),
    .io_sortedFrequency_15(sort_io_sortedFrequency_15),
    .io_sortedFrequency_16(sort_io_sortedFrequency_16),
    .io_sortedFrequency_17(sort_io_sortedFrequency_17),
    .io_sortedFrequency_18(sort_io_sortedFrequency_18),
    .io_sortedFrequency_19(sort_io_sortedFrequency_19),
    .io_sortedFrequency_20(sort_io_sortedFrequency_20),
    .io_sortedFrequency_21(sort_io_sortedFrequency_21),
    .io_sortedFrequency_22(sort_io_sortedFrequency_22),
    .io_sortedFrequency_23(sort_io_sortedFrequency_23),
    .io_sortedFrequency_24(sort_io_sortedFrequency_24),
    .io_sortedFrequency_25(sort_io_sortedFrequency_25),
    .io_sortedFrequency_26(sort_io_sortedFrequency_26),
    .io_sortedFrequency_27(sort_io_sortedFrequency_27),
    .io_sortedFrequency_28(sort_io_sortedFrequency_28),
    .io_sortedFrequency_29(sort_io_sortedFrequency_29),
    .io_sortedFrequency_30(sort_io_sortedFrequency_30),
    .io_sortedFrequency_31(sort_io_sortedFrequency_31),
    .io_sortedCharacter_0(sort_io_sortedCharacter_0),
    .io_sortedCharacter_1(sort_io_sortedCharacter_1),
    .io_sortedCharacter_2(sort_io_sortedCharacter_2),
    .io_sortedCharacter_3(sort_io_sortedCharacter_3),
    .io_sortedCharacter_4(sort_io_sortedCharacter_4),
    .io_sortedCharacter_5(sort_io_sortedCharacter_5),
    .io_sortedCharacter_6(sort_io_sortedCharacter_6),
    .io_sortedCharacter_7(sort_io_sortedCharacter_7),
    .io_sortedCharacter_8(sort_io_sortedCharacter_8),
    .io_sortedCharacter_9(sort_io_sortedCharacter_9),
    .io_sortedCharacter_10(sort_io_sortedCharacter_10),
    .io_sortedCharacter_11(sort_io_sortedCharacter_11),
    .io_sortedCharacter_12(sort_io_sortedCharacter_12),
    .io_sortedCharacter_13(sort_io_sortedCharacter_13),
    .io_sortedCharacter_14(sort_io_sortedCharacter_14),
    .io_sortedCharacter_15(sort_io_sortedCharacter_15),
    .io_sortedCharacter_16(sort_io_sortedCharacter_16),
    .io_sortedCharacter_17(sort_io_sortedCharacter_17),
    .io_sortedCharacter_18(sort_io_sortedCharacter_18),
    .io_sortedCharacter_19(sort_io_sortedCharacter_19),
    .io_sortedCharacter_20(sort_io_sortedCharacter_20),
    .io_sortedCharacter_21(sort_io_sortedCharacter_21),
    .io_sortedCharacter_22(sort_io_sortedCharacter_22),
    .io_sortedCharacter_23(sort_io_sortedCharacter_23),
    .io_sortedCharacter_24(sort_io_sortedCharacter_24),
    .io_sortedCharacter_25(sort_io_sortedCharacter_25),
    .io_sortedCharacter_26(sort_io_sortedCharacter_26),
    .io_sortedCharacter_27(sort_io_sortedCharacter_27),
    .io_sortedCharacter_28(sort_io_sortedCharacter_28),
    .io_sortedCharacter_29(sort_io_sortedCharacter_29),
    .io_sortedCharacter_30(sort_io_sortedCharacter_30),
    .io_sortedCharacter_31(sort_io_sortedCharacter_31),
    .io_finished(sort_io_finished)
  );
  assign io_input_currentByteOut = input__io_input_currentByteOut; // @[characterFrequencyModule.scala 42:18]
  assign io_input_ready = input__io_input_ready; // @[characterFrequencyModule.scala 42:18]
  assign io_outputs_sortedFrequency_0 = sort_io_sortedFrequency_0; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_1 = sort_io_sortedFrequency_1; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_2 = sort_io_sortedFrequency_2; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_3 = sort_io_sortedFrequency_3; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_4 = sort_io_sortedFrequency_4; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_5 = sort_io_sortedFrequency_5; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_6 = sort_io_sortedFrequency_6; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_7 = sort_io_sortedFrequency_7; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_8 = sort_io_sortedFrequency_8; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_9 = sort_io_sortedFrequency_9; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_10 = sort_io_sortedFrequency_10; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_11 = sort_io_sortedFrequency_11; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_12 = sort_io_sortedFrequency_12; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_13 = sort_io_sortedFrequency_13; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_14 = sort_io_sortedFrequency_14; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_15 = sort_io_sortedFrequency_15; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_16 = sort_io_sortedFrequency_16; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_17 = sort_io_sortedFrequency_17; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_18 = sort_io_sortedFrequency_18; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_19 = sort_io_sortedFrequency_19; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_20 = sort_io_sortedFrequency_20; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_21 = sort_io_sortedFrequency_21; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_22 = sort_io_sortedFrequency_22; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_23 = sort_io_sortedFrequency_23; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_24 = sort_io_sortedFrequency_24; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_25 = sort_io_sortedFrequency_25; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_26 = sort_io_sortedFrequency_26; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_27 = sort_io_sortedFrequency_27; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_28 = sort_io_sortedFrequency_28; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_29 = sort_io_sortedFrequency_29; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_30 = sort_io_sortedFrequency_30; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedFrequency_31 = sort_io_sortedFrequency_31; // @[characterFrequencyModule.scala 46:30]
  assign io_outputs_sortedCharacter_0 = sort_io_sortedCharacter_0; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_1 = sort_io_sortedCharacter_1; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_2 = sort_io_sortedCharacter_2; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_3 = sort_io_sortedCharacter_3; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_4 = sort_io_sortedCharacter_4; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_5 = sort_io_sortedCharacter_5; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_6 = sort_io_sortedCharacter_6; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_7 = sort_io_sortedCharacter_7; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_8 = sort_io_sortedCharacter_8; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_9 = sort_io_sortedCharacter_9; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_10 = sort_io_sortedCharacter_10; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_11 = sort_io_sortedCharacter_11; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_12 = sort_io_sortedCharacter_12; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_13 = sort_io_sortedCharacter_13; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_14 = sort_io_sortedCharacter_14; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_15 = sort_io_sortedCharacter_15; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_16 = sort_io_sortedCharacter_16; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_17 = sort_io_sortedCharacter_17; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_18 = sort_io_sortedCharacter_18; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_19 = sort_io_sortedCharacter_19; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_20 = sort_io_sortedCharacter_20; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_21 = sort_io_sortedCharacter_21; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_22 = sort_io_sortedCharacter_22; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_23 = sort_io_sortedCharacter_23; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_24 = sort_io_sortedCharacter_24; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_25 = sort_io_sortedCharacter_25; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_26 = sort_io_sortedCharacter_26; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_27 = sort_io_sortedCharacter_27; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_28 = sort_io_sortedCharacter_28; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_29 = sort_io_sortedCharacter_29; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_30 = sort_io_sortedCharacter_30; // @[characterFrequencyModule.scala 47:30]
  assign io_outputs_sortedCharacter_31 = sort_io_sortedCharacter_31; // @[characterFrequencyModule.scala 47:30]
  assign io_finished = sort_io_finished; // @[characterFrequencyModule.scala 39:15]
  assign input__io_input_dataIn_0 = io_input_dataIn_0; // @[characterFrequencyModule.scala 42:18]
  assign input__io_input_valid = io_input_valid; // @[characterFrequencyModule.scala 42:18]
  assign input__io_currentByte = count_io_currentByte; // @[characterFrequencyModule.scala 45:24]
  assign input__io_dataOut_ready = count_io_dataIn_ready; // @[characterFrequencyModule.scala 41:19]
  assign count_clock = clock;
  assign count_reset = reset;
  assign count_io_start = io_start; // @[characterFrequencyModule.scala 44:18]
  assign count_io_dataIn_bits_0 = input__io_dataOut_bits_0; // @[characterFrequencyModule.scala 41:19]
  assign sort_clock = clock;
  assign sort_reset = reset;
  assign sort_io_start = count_io_finished & _T; // @[characterFrequencyModule.scala 38:17]
  assign sort_io_dataIn_0 = count_io_frequencies_0; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_1 = count_io_frequencies_1; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_2 = count_io_frequencies_2; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_3 = count_io_frequencies_3; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_4 = count_io_frequencies_4; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_5 = count_io_frequencies_5; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_6 = count_io_frequencies_6; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_7 = count_io_frequencies_7; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_8 = count_io_frequencies_8; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_9 = count_io_frequencies_9; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_10 = count_io_frequencies_10; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_11 = count_io_frequencies_11; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_12 = count_io_frequencies_12; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_13 = count_io_frequencies_13; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_14 = count_io_frequencies_14; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_15 = count_io_frequencies_15; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_16 = count_io_frequencies_16; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_17 = count_io_frequencies_17; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_18 = count_io_frequencies_18; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_19 = count_io_frequencies_19; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_20 = count_io_frequencies_20; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_21 = count_io_frequencies_21; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_22 = count_io_frequencies_22; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_23 = count_io_frequencies_23; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_24 = count_io_frequencies_24; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_25 = count_io_frequencies_25; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_26 = count_io_frequencies_26; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_27 = count_io_frequencies_27; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_28 = count_io_frequencies_28; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_29 = count_io_frequencies_29; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_30 = count_io_frequencies_30; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_31 = count_io_frequencies_31; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_32 = count_io_frequencies_32; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_33 = count_io_frequencies_33; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_34 = count_io_frequencies_34; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_35 = count_io_frequencies_35; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_36 = count_io_frequencies_36; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_37 = count_io_frequencies_37; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_38 = count_io_frequencies_38; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_39 = count_io_frequencies_39; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_40 = count_io_frequencies_40; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_41 = count_io_frequencies_41; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_42 = count_io_frequencies_42; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_43 = count_io_frequencies_43; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_44 = count_io_frequencies_44; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_45 = count_io_frequencies_45; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_46 = count_io_frequencies_46; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_47 = count_io_frequencies_47; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_48 = count_io_frequencies_48; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_49 = count_io_frequencies_49; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_50 = count_io_frequencies_50; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_51 = count_io_frequencies_51; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_52 = count_io_frequencies_52; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_53 = count_io_frequencies_53; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_54 = count_io_frequencies_54; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_55 = count_io_frequencies_55; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_56 = count_io_frequencies_56; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_57 = count_io_frequencies_57; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_58 = count_io_frequencies_58; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_59 = count_io_frequencies_59; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_60 = count_io_frequencies_60; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_61 = count_io_frequencies_61; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_62 = count_io_frequencies_62; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_63 = count_io_frequencies_63; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_64 = count_io_frequencies_64; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_65 = count_io_frequencies_65; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_66 = count_io_frequencies_66; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_67 = count_io_frequencies_67; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_68 = count_io_frequencies_68; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_69 = count_io_frequencies_69; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_70 = count_io_frequencies_70; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_71 = count_io_frequencies_71; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_72 = count_io_frequencies_72; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_73 = count_io_frequencies_73; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_74 = count_io_frequencies_74; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_75 = count_io_frequencies_75; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_76 = count_io_frequencies_76; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_77 = count_io_frequencies_77; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_78 = count_io_frequencies_78; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_79 = count_io_frequencies_79; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_80 = count_io_frequencies_80; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_81 = count_io_frequencies_81; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_82 = count_io_frequencies_82; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_83 = count_io_frequencies_83; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_84 = count_io_frequencies_84; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_85 = count_io_frequencies_85; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_86 = count_io_frequencies_86; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_87 = count_io_frequencies_87; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_88 = count_io_frequencies_88; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_89 = count_io_frequencies_89; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_90 = count_io_frequencies_90; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_91 = count_io_frequencies_91; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_92 = count_io_frequencies_92; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_93 = count_io_frequencies_93; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_94 = count_io_frequencies_94; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_95 = count_io_frequencies_95; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_96 = count_io_frequencies_96; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_97 = count_io_frequencies_97; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_98 = count_io_frequencies_98; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_99 = count_io_frequencies_99; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_100 = count_io_frequencies_100; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_101 = count_io_frequencies_101; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_102 = count_io_frequencies_102; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_103 = count_io_frequencies_103; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_104 = count_io_frequencies_104; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_105 = count_io_frequencies_105; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_106 = count_io_frequencies_106; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_107 = count_io_frequencies_107; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_108 = count_io_frequencies_108; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_109 = count_io_frequencies_109; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_110 = count_io_frequencies_110; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_111 = count_io_frequencies_111; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_112 = count_io_frequencies_112; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_113 = count_io_frequencies_113; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_114 = count_io_frequencies_114; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_115 = count_io_frequencies_115; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_116 = count_io_frequencies_116; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_117 = count_io_frequencies_117; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_118 = count_io_frequencies_118; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_119 = count_io_frequencies_119; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_120 = count_io_frequencies_120; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_121 = count_io_frequencies_121; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_122 = count_io_frequencies_122; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_123 = count_io_frequencies_123; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_124 = count_io_frequencies_124; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_125 = count_io_frequencies_125; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_126 = count_io_frequencies_126; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_127 = count_io_frequencies_127; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_128 = count_io_frequencies_128; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_129 = count_io_frequencies_129; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_130 = count_io_frequencies_130; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_131 = count_io_frequencies_131; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_132 = count_io_frequencies_132; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_133 = count_io_frequencies_133; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_134 = count_io_frequencies_134; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_135 = count_io_frequencies_135; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_136 = count_io_frequencies_136; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_137 = count_io_frequencies_137; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_138 = count_io_frequencies_138; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_139 = count_io_frequencies_139; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_140 = count_io_frequencies_140; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_141 = count_io_frequencies_141; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_142 = count_io_frequencies_142; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_143 = count_io_frequencies_143; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_144 = count_io_frequencies_144; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_145 = count_io_frequencies_145; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_146 = count_io_frequencies_146; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_147 = count_io_frequencies_147; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_148 = count_io_frequencies_148; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_149 = count_io_frequencies_149; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_150 = count_io_frequencies_150; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_151 = count_io_frequencies_151; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_152 = count_io_frequencies_152; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_153 = count_io_frequencies_153; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_154 = count_io_frequencies_154; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_155 = count_io_frequencies_155; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_156 = count_io_frequencies_156; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_157 = count_io_frequencies_157; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_158 = count_io_frequencies_158; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_159 = count_io_frequencies_159; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_160 = count_io_frequencies_160; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_161 = count_io_frequencies_161; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_162 = count_io_frequencies_162; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_163 = count_io_frequencies_163; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_164 = count_io_frequencies_164; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_165 = count_io_frequencies_165; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_166 = count_io_frequencies_166; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_167 = count_io_frequencies_167; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_168 = count_io_frequencies_168; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_169 = count_io_frequencies_169; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_170 = count_io_frequencies_170; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_171 = count_io_frequencies_171; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_172 = count_io_frequencies_172; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_173 = count_io_frequencies_173; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_174 = count_io_frequencies_174; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_175 = count_io_frequencies_175; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_176 = count_io_frequencies_176; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_177 = count_io_frequencies_177; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_178 = count_io_frequencies_178; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_179 = count_io_frequencies_179; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_180 = count_io_frequencies_180; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_181 = count_io_frequencies_181; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_182 = count_io_frequencies_182; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_183 = count_io_frequencies_183; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_184 = count_io_frequencies_184; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_185 = count_io_frequencies_185; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_186 = count_io_frequencies_186; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_187 = count_io_frequencies_187; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_188 = count_io_frequencies_188; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_189 = count_io_frequencies_189; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_190 = count_io_frequencies_190; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_191 = count_io_frequencies_191; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_192 = count_io_frequencies_192; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_193 = count_io_frequencies_193; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_194 = count_io_frequencies_194; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_195 = count_io_frequencies_195; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_196 = count_io_frequencies_196; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_197 = count_io_frequencies_197; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_198 = count_io_frequencies_198; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_199 = count_io_frequencies_199; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_200 = count_io_frequencies_200; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_201 = count_io_frequencies_201; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_202 = count_io_frequencies_202; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_203 = count_io_frequencies_203; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_204 = count_io_frequencies_204; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_205 = count_io_frequencies_205; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_206 = count_io_frequencies_206; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_207 = count_io_frequencies_207; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_208 = count_io_frequencies_208; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_209 = count_io_frequencies_209; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_210 = count_io_frequencies_210; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_211 = count_io_frequencies_211; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_212 = count_io_frequencies_212; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_213 = count_io_frequencies_213; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_214 = count_io_frequencies_214; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_215 = count_io_frequencies_215; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_216 = count_io_frequencies_216; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_217 = count_io_frequencies_217; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_218 = count_io_frequencies_218; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_219 = count_io_frequencies_219; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_220 = count_io_frequencies_220; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_221 = count_io_frequencies_221; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_222 = count_io_frequencies_222; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_223 = count_io_frequencies_223; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_224 = count_io_frequencies_224; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_225 = count_io_frequencies_225; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_226 = count_io_frequencies_226; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_227 = count_io_frequencies_227; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_228 = count_io_frequencies_228; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_229 = count_io_frequencies_229; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_230 = count_io_frequencies_230; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_231 = count_io_frequencies_231; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_232 = count_io_frequencies_232; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_233 = count_io_frequencies_233; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_234 = count_io_frequencies_234; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_235 = count_io_frequencies_235; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_236 = count_io_frequencies_236; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_237 = count_io_frequencies_237; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_238 = count_io_frequencies_238; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_239 = count_io_frequencies_239; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_240 = count_io_frequencies_240; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_241 = count_io_frequencies_241; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_242 = count_io_frequencies_242; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_243 = count_io_frequencies_243; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_244 = count_io_frequencies_244; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_245 = count_io_frequencies_245; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_246 = count_io_frequencies_246; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_247 = count_io_frequencies_247; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_248 = count_io_frequencies_248; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_249 = count_io_frequencies_249; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_250 = count_io_frequencies_250; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_251 = count_io_frequencies_251; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_252 = count_io_frequencies_252; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_253 = count_io_frequencies_253; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_254 = count_io_frequencies_254; // @[characterFrequencyModule.scala 40:18]
  assign sort_io_dataIn_255 = count_io_frequencies_255; // @[characterFrequencyModule.scala 40:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  previousCountFinished = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    previousCountFinished <= count_io_finished;
  end
endmodule
module treeGenerator(
  input         clock,
  input         reset,
  input         io_start,
  input  [12:0] io_inputs_sortedFrequency_0,
  input  [12:0] io_inputs_sortedFrequency_1,
  input  [12:0] io_inputs_sortedFrequency_2,
  input  [12:0] io_inputs_sortedFrequency_3,
  input  [12:0] io_inputs_sortedFrequency_4,
  input  [12:0] io_inputs_sortedFrequency_5,
  input  [12:0] io_inputs_sortedFrequency_6,
  input  [12:0] io_inputs_sortedFrequency_7,
  input  [12:0] io_inputs_sortedFrequency_8,
  input  [12:0] io_inputs_sortedFrequency_9,
  input  [12:0] io_inputs_sortedFrequency_10,
  input  [12:0] io_inputs_sortedFrequency_11,
  input  [12:0] io_inputs_sortedFrequency_12,
  input  [12:0] io_inputs_sortedFrequency_13,
  input  [12:0] io_inputs_sortedFrequency_14,
  input  [12:0] io_inputs_sortedFrequency_15,
  input  [12:0] io_inputs_sortedFrequency_16,
  input  [12:0] io_inputs_sortedFrequency_17,
  input  [12:0] io_inputs_sortedFrequency_18,
  input  [12:0] io_inputs_sortedFrequency_19,
  input  [12:0] io_inputs_sortedFrequency_20,
  input  [12:0] io_inputs_sortedFrequency_21,
  input  [12:0] io_inputs_sortedFrequency_22,
  input  [12:0] io_inputs_sortedFrequency_23,
  input  [12:0] io_inputs_sortedFrequency_24,
  input  [12:0] io_inputs_sortedFrequency_25,
  input  [12:0] io_inputs_sortedFrequency_26,
  input  [12:0] io_inputs_sortedFrequency_27,
  input  [12:0] io_inputs_sortedFrequency_28,
  input  [12:0] io_inputs_sortedFrequency_29,
  input  [12:0] io_inputs_sortedFrequency_30,
  input  [12:0] io_inputs_sortedFrequency_31,
  input  [8:0]  io_inputs_sortedCharacter_0,
  input  [8:0]  io_inputs_sortedCharacter_1,
  input  [8:0]  io_inputs_sortedCharacter_2,
  input  [8:0]  io_inputs_sortedCharacter_3,
  input  [8:0]  io_inputs_sortedCharacter_4,
  input  [8:0]  io_inputs_sortedCharacter_5,
  input  [8:0]  io_inputs_sortedCharacter_6,
  input  [8:0]  io_inputs_sortedCharacter_7,
  input  [8:0]  io_inputs_sortedCharacter_8,
  input  [8:0]  io_inputs_sortedCharacter_9,
  input  [8:0]  io_inputs_sortedCharacter_10,
  input  [8:0]  io_inputs_sortedCharacter_11,
  input  [8:0]  io_inputs_sortedCharacter_12,
  input  [8:0]  io_inputs_sortedCharacter_13,
  input  [8:0]  io_inputs_sortedCharacter_14,
  input  [8:0]  io_inputs_sortedCharacter_15,
  input  [8:0]  io_inputs_sortedCharacter_16,
  input  [8:0]  io_inputs_sortedCharacter_17,
  input  [8:0]  io_inputs_sortedCharacter_18,
  input  [8:0]  io_inputs_sortedCharacter_19,
  input  [8:0]  io_inputs_sortedCharacter_20,
  input  [8:0]  io_inputs_sortedCharacter_21,
  input  [8:0]  io_inputs_sortedCharacter_22,
  input  [8:0]  io_inputs_sortedCharacter_23,
  input  [8:0]  io_inputs_sortedCharacter_24,
  input  [8:0]  io_inputs_sortedCharacter_25,
  input  [8:0]  io_inputs_sortedCharacter_26,
  input  [8:0]  io_inputs_sortedCharacter_27,
  input  [8:0]  io_inputs_sortedCharacter_28,
  input  [8:0]  io_inputs_sortedCharacter_29,
  input  [8:0]  io_inputs_sortedCharacter_30,
  input  [8:0]  io_inputs_sortedCharacter_31,
  output [8:0]  io_outputs_leftNode_0,
  output [8:0]  io_outputs_leftNode_1,
  output [8:0]  io_outputs_leftNode_2,
  output [8:0]  io_outputs_leftNode_3,
  output [8:0]  io_outputs_leftNode_4,
  output [8:0]  io_outputs_leftNode_5,
  output [8:0]  io_outputs_leftNode_6,
  output [8:0]  io_outputs_leftNode_7,
  output [8:0]  io_outputs_leftNode_8,
  output [8:0]  io_outputs_leftNode_9,
  output [8:0]  io_outputs_leftNode_10,
  output [8:0]  io_outputs_leftNode_11,
  output [8:0]  io_outputs_leftNode_12,
  output [8:0]  io_outputs_leftNode_13,
  output [8:0]  io_outputs_leftNode_14,
  output [8:0]  io_outputs_leftNode_15,
  output [8:0]  io_outputs_leftNode_16,
  output [8:0]  io_outputs_leftNode_17,
  output [8:0]  io_outputs_leftNode_18,
  output [8:0]  io_outputs_leftNode_19,
  output [8:0]  io_outputs_leftNode_20,
  output [8:0]  io_outputs_leftNode_21,
  output [8:0]  io_outputs_leftNode_22,
  output [8:0]  io_outputs_leftNode_23,
  output [8:0]  io_outputs_leftNode_24,
  output [8:0]  io_outputs_leftNode_25,
  output [8:0]  io_outputs_leftNode_26,
  output [8:0]  io_outputs_leftNode_27,
  output [8:0]  io_outputs_leftNode_28,
  output [8:0]  io_outputs_leftNode_29,
  output [8:0]  io_outputs_leftNode_30,
  output [8:0]  io_outputs_leftNode_31,
  output [8:0]  io_outputs_leftNode_32,
  output [8:0]  io_outputs_leftNode_33,
  output [8:0]  io_outputs_leftNode_34,
  output [8:0]  io_outputs_leftNode_35,
  output [8:0]  io_outputs_leftNode_36,
  output [8:0]  io_outputs_leftNode_37,
  output [8:0]  io_outputs_leftNode_38,
  output [8:0]  io_outputs_leftNode_39,
  output [8:0]  io_outputs_leftNode_40,
  output [8:0]  io_outputs_leftNode_41,
  output [8:0]  io_outputs_leftNode_42,
  output [8:0]  io_outputs_leftNode_43,
  output [8:0]  io_outputs_leftNode_44,
  output [8:0]  io_outputs_leftNode_45,
  output [8:0]  io_outputs_leftNode_46,
  output [8:0]  io_outputs_leftNode_47,
  output [8:0]  io_outputs_leftNode_48,
  output [8:0]  io_outputs_leftNode_49,
  output [8:0]  io_outputs_leftNode_50,
  output [8:0]  io_outputs_leftNode_51,
  output [8:0]  io_outputs_leftNode_52,
  output [8:0]  io_outputs_leftNode_53,
  output [8:0]  io_outputs_leftNode_54,
  output [8:0]  io_outputs_leftNode_55,
  output [8:0]  io_outputs_leftNode_56,
  output [8:0]  io_outputs_leftNode_57,
  output [8:0]  io_outputs_leftNode_58,
  output [8:0]  io_outputs_leftNode_59,
  output [8:0]  io_outputs_leftNode_60,
  output [8:0]  io_outputs_leftNode_61,
  output [8:0]  io_outputs_leftNode_62,
  output [8:0]  io_outputs_leftNode_63,
  output [8:0]  io_outputs_rightNode_0,
  output [8:0]  io_outputs_rightNode_1,
  output [8:0]  io_outputs_rightNode_2,
  output [8:0]  io_outputs_rightNode_3,
  output [8:0]  io_outputs_rightNode_4,
  output [8:0]  io_outputs_rightNode_5,
  output [8:0]  io_outputs_rightNode_6,
  output [8:0]  io_outputs_rightNode_7,
  output [8:0]  io_outputs_rightNode_8,
  output [8:0]  io_outputs_rightNode_9,
  output [8:0]  io_outputs_rightNode_10,
  output [8:0]  io_outputs_rightNode_11,
  output [8:0]  io_outputs_rightNode_12,
  output [8:0]  io_outputs_rightNode_13,
  output [8:0]  io_outputs_rightNode_14,
  output [8:0]  io_outputs_rightNode_15,
  output [8:0]  io_outputs_rightNode_16,
  output [8:0]  io_outputs_rightNode_17,
  output [8:0]  io_outputs_rightNode_18,
  output [8:0]  io_outputs_rightNode_19,
  output [8:0]  io_outputs_rightNode_20,
  output [8:0]  io_outputs_rightNode_21,
  output [8:0]  io_outputs_rightNode_22,
  output [8:0]  io_outputs_rightNode_23,
  output [8:0]  io_outputs_rightNode_24,
  output [8:0]  io_outputs_rightNode_25,
  output [8:0]  io_outputs_rightNode_26,
  output [8:0]  io_outputs_rightNode_27,
  output [8:0]  io_outputs_rightNode_28,
  output [8:0]  io_outputs_rightNode_29,
  output [8:0]  io_outputs_rightNode_30,
  output [8:0]  io_outputs_rightNode_31,
  output [8:0]  io_outputs_rightNode_32,
  output [8:0]  io_outputs_rightNode_33,
  output [8:0]  io_outputs_rightNode_34,
  output [8:0]  io_outputs_rightNode_35,
  output [8:0]  io_outputs_rightNode_36,
  output [8:0]  io_outputs_rightNode_37,
  output [8:0]  io_outputs_rightNode_38,
  output [8:0]  io_outputs_rightNode_39,
  output [8:0]  io_outputs_rightNode_40,
  output [8:0]  io_outputs_rightNode_41,
  output [8:0]  io_outputs_rightNode_42,
  output [8:0]  io_outputs_rightNode_43,
  output [8:0]  io_outputs_rightNode_44,
  output [8:0]  io_outputs_rightNode_45,
  output [8:0]  io_outputs_rightNode_46,
  output [8:0]  io_outputs_rightNode_47,
  output [8:0]  io_outputs_rightNode_48,
  output [8:0]  io_outputs_rightNode_49,
  output [8:0]  io_outputs_rightNode_50,
  output [8:0]  io_outputs_rightNode_51,
  output [8:0]  io_outputs_rightNode_52,
  output [8:0]  io_outputs_rightNode_53,
  output [8:0]  io_outputs_rightNode_54,
  output [8:0]  io_outputs_rightNode_55,
  output [8:0]  io_outputs_rightNode_56,
  output [8:0]  io_outputs_rightNode_57,
  output [8:0]  io_outputs_rightNode_58,
  output [8:0]  io_outputs_rightNode_59,
  output [8:0]  io_outputs_rightNode_60,
  output [8:0]  io_outputs_rightNode_61,
  output [8:0]  io_outputs_rightNode_62,
  output [8:0]  io_outputs_rightNode_63,
  output        io_outputs_leftNodeIsCharacter_0,
  output        io_outputs_leftNodeIsCharacter_1,
  output        io_outputs_leftNodeIsCharacter_2,
  output        io_outputs_leftNodeIsCharacter_3,
  output        io_outputs_leftNodeIsCharacter_4,
  output        io_outputs_leftNodeIsCharacter_5,
  output        io_outputs_leftNodeIsCharacter_6,
  output        io_outputs_leftNodeIsCharacter_7,
  output        io_outputs_leftNodeIsCharacter_8,
  output        io_outputs_leftNodeIsCharacter_9,
  output        io_outputs_leftNodeIsCharacter_10,
  output        io_outputs_leftNodeIsCharacter_11,
  output        io_outputs_leftNodeIsCharacter_12,
  output        io_outputs_leftNodeIsCharacter_13,
  output        io_outputs_leftNodeIsCharacter_14,
  output        io_outputs_leftNodeIsCharacter_15,
  output        io_outputs_leftNodeIsCharacter_16,
  output        io_outputs_leftNodeIsCharacter_17,
  output        io_outputs_leftNodeIsCharacter_18,
  output        io_outputs_leftNodeIsCharacter_19,
  output        io_outputs_leftNodeIsCharacter_20,
  output        io_outputs_leftNodeIsCharacter_21,
  output        io_outputs_leftNodeIsCharacter_22,
  output        io_outputs_leftNodeIsCharacter_23,
  output        io_outputs_leftNodeIsCharacter_24,
  output        io_outputs_leftNodeIsCharacter_25,
  output        io_outputs_leftNodeIsCharacter_26,
  output        io_outputs_leftNodeIsCharacter_27,
  output        io_outputs_leftNodeIsCharacter_28,
  output        io_outputs_leftNodeIsCharacter_29,
  output        io_outputs_leftNodeIsCharacter_30,
  output        io_outputs_leftNodeIsCharacter_31,
  output        io_outputs_leftNodeIsCharacter_32,
  output        io_outputs_leftNodeIsCharacter_33,
  output        io_outputs_leftNodeIsCharacter_34,
  output        io_outputs_leftNodeIsCharacter_35,
  output        io_outputs_leftNodeIsCharacter_36,
  output        io_outputs_leftNodeIsCharacter_37,
  output        io_outputs_leftNodeIsCharacter_38,
  output        io_outputs_leftNodeIsCharacter_39,
  output        io_outputs_leftNodeIsCharacter_40,
  output        io_outputs_leftNodeIsCharacter_41,
  output        io_outputs_leftNodeIsCharacter_42,
  output        io_outputs_leftNodeIsCharacter_43,
  output        io_outputs_leftNodeIsCharacter_44,
  output        io_outputs_leftNodeIsCharacter_45,
  output        io_outputs_leftNodeIsCharacter_46,
  output        io_outputs_leftNodeIsCharacter_47,
  output        io_outputs_leftNodeIsCharacter_48,
  output        io_outputs_leftNodeIsCharacter_49,
  output        io_outputs_leftNodeIsCharacter_50,
  output        io_outputs_leftNodeIsCharacter_51,
  output        io_outputs_leftNodeIsCharacter_52,
  output        io_outputs_leftNodeIsCharacter_53,
  output        io_outputs_leftNodeIsCharacter_54,
  output        io_outputs_leftNodeIsCharacter_55,
  output        io_outputs_leftNodeIsCharacter_56,
  output        io_outputs_leftNodeIsCharacter_57,
  output        io_outputs_leftNodeIsCharacter_58,
  output        io_outputs_leftNodeIsCharacter_59,
  output        io_outputs_leftNodeIsCharacter_60,
  output        io_outputs_leftNodeIsCharacter_61,
  output        io_outputs_leftNodeIsCharacter_62,
  output        io_outputs_leftNodeIsCharacter_63,
  output        io_outputs_rightNodeIsCharacter_0,
  output        io_outputs_rightNodeIsCharacter_1,
  output        io_outputs_rightNodeIsCharacter_2,
  output        io_outputs_rightNodeIsCharacter_3,
  output        io_outputs_rightNodeIsCharacter_4,
  output        io_outputs_rightNodeIsCharacter_5,
  output        io_outputs_rightNodeIsCharacter_6,
  output        io_outputs_rightNodeIsCharacter_7,
  output        io_outputs_rightNodeIsCharacter_8,
  output        io_outputs_rightNodeIsCharacter_9,
  output        io_outputs_rightNodeIsCharacter_10,
  output        io_outputs_rightNodeIsCharacter_11,
  output        io_outputs_rightNodeIsCharacter_12,
  output        io_outputs_rightNodeIsCharacter_13,
  output        io_outputs_rightNodeIsCharacter_14,
  output        io_outputs_rightNodeIsCharacter_15,
  output        io_outputs_rightNodeIsCharacter_16,
  output        io_outputs_rightNodeIsCharacter_17,
  output        io_outputs_rightNodeIsCharacter_18,
  output        io_outputs_rightNodeIsCharacter_19,
  output        io_outputs_rightNodeIsCharacter_20,
  output        io_outputs_rightNodeIsCharacter_21,
  output        io_outputs_rightNodeIsCharacter_22,
  output        io_outputs_rightNodeIsCharacter_23,
  output        io_outputs_rightNodeIsCharacter_24,
  output        io_outputs_rightNodeIsCharacter_25,
  output        io_outputs_rightNodeIsCharacter_26,
  output        io_outputs_rightNodeIsCharacter_27,
  output        io_outputs_rightNodeIsCharacter_28,
  output        io_outputs_rightNodeIsCharacter_29,
  output        io_outputs_rightNodeIsCharacter_30,
  output        io_outputs_rightNodeIsCharacter_31,
  output        io_outputs_rightNodeIsCharacter_32,
  output        io_outputs_rightNodeIsCharacter_33,
  output        io_outputs_rightNodeIsCharacter_34,
  output        io_outputs_rightNodeIsCharacter_35,
  output        io_outputs_rightNodeIsCharacter_36,
  output        io_outputs_rightNodeIsCharacter_37,
  output        io_outputs_rightNodeIsCharacter_38,
  output        io_outputs_rightNodeIsCharacter_39,
  output        io_outputs_rightNodeIsCharacter_40,
  output        io_outputs_rightNodeIsCharacter_41,
  output        io_outputs_rightNodeIsCharacter_42,
  output        io_outputs_rightNodeIsCharacter_43,
  output        io_outputs_rightNodeIsCharacter_44,
  output        io_outputs_rightNodeIsCharacter_45,
  output        io_outputs_rightNodeIsCharacter_46,
  output        io_outputs_rightNodeIsCharacter_47,
  output        io_outputs_rightNodeIsCharacter_48,
  output        io_outputs_rightNodeIsCharacter_49,
  output        io_outputs_rightNodeIsCharacter_50,
  output        io_outputs_rightNodeIsCharacter_51,
  output        io_outputs_rightNodeIsCharacter_52,
  output        io_outputs_rightNodeIsCharacter_53,
  output        io_outputs_rightNodeIsCharacter_54,
  output        io_outputs_rightNodeIsCharacter_55,
  output        io_outputs_rightNodeIsCharacter_56,
  output        io_outputs_rightNodeIsCharacter_57,
  output        io_outputs_rightNodeIsCharacter_58,
  output        io_outputs_rightNodeIsCharacter_59,
  output        io_outputs_rightNodeIsCharacter_60,
  output        io_outputs_rightNodeIsCharacter_61,
  output        io_outputs_rightNodeIsCharacter_62,
  output        io_outputs_rightNodeIsCharacter_63,
  output [6:0]  io_outputs_validNodes,
  output [5:0]  io_outputs_validCharacters,
  output        io_finished
);
  reg [12:0] frequency_0; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_0;
  reg [12:0] frequency_1; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_1;
  reg [12:0] frequency_2; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_2;
  reg [12:0] frequency_3; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_3;
  reg [12:0] frequency_4; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_4;
  reg [12:0] frequency_5; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_5;
  reg [12:0] frequency_6; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_6;
  reg [12:0] frequency_7; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_7;
  reg [12:0] frequency_8; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_8;
  reg [12:0] frequency_9; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_9;
  reg [12:0] frequency_10; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_10;
  reg [12:0] frequency_11; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_11;
  reg [12:0] frequency_12; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_12;
  reg [12:0] frequency_13; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_13;
  reg [12:0] frequency_14; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_14;
  reg [12:0] frequency_15; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_15;
  reg [12:0] frequency_16; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_16;
  reg [12:0] frequency_17; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_17;
  reg [12:0] frequency_18; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_18;
  reg [12:0] frequency_19; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_19;
  reg [12:0] frequency_20; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_20;
  reg [12:0] frequency_21; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_21;
  reg [12:0] frequency_22; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_22;
  reg [12:0] frequency_23; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_23;
  reg [12:0] frequency_24; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_24;
  reg [12:0] frequency_25; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_25;
  reg [12:0] frequency_26; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_26;
  reg [12:0] frequency_27; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_27;
  reg [12:0] frequency_28; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_28;
  reg [12:0] frequency_29; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_29;
  reg [12:0] frequency_30; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_30;
  reg [12:0] frequency_31; // @[treeGenerator.scala 22:22]
  reg [31:0] _RAND_31;
  reg [8:0] pointerOrCharacter_0; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_32;
  reg [8:0] pointerOrCharacter_1; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_33;
  reg [8:0] pointerOrCharacter_2; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_34;
  reg [8:0] pointerOrCharacter_3; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_35;
  reg [8:0] pointerOrCharacter_4; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_36;
  reg [8:0] pointerOrCharacter_5; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_37;
  reg [8:0] pointerOrCharacter_6; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_38;
  reg [8:0] pointerOrCharacter_7; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_39;
  reg [8:0] pointerOrCharacter_8; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_40;
  reg [8:0] pointerOrCharacter_9; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_41;
  reg [8:0] pointerOrCharacter_10; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_42;
  reg [8:0] pointerOrCharacter_11; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_43;
  reg [8:0] pointerOrCharacter_12; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_44;
  reg [8:0] pointerOrCharacter_13; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_45;
  reg [8:0] pointerOrCharacter_14; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_46;
  reg [8:0] pointerOrCharacter_15; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_47;
  reg [8:0] pointerOrCharacter_16; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_48;
  reg [8:0] pointerOrCharacter_17; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_49;
  reg [8:0] pointerOrCharacter_18; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_50;
  reg [8:0] pointerOrCharacter_19; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_51;
  reg [8:0] pointerOrCharacter_20; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_52;
  reg [8:0] pointerOrCharacter_21; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_53;
  reg [8:0] pointerOrCharacter_22; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_54;
  reg [8:0] pointerOrCharacter_23; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_55;
  reg [8:0] pointerOrCharacter_24; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_56;
  reg [8:0] pointerOrCharacter_25; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_57;
  reg [8:0] pointerOrCharacter_26; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_58;
  reg [8:0] pointerOrCharacter_27; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_59;
  reg [8:0] pointerOrCharacter_28; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_60;
  reg [8:0] pointerOrCharacter_29; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_61;
  reg [8:0] pointerOrCharacter_30; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_62;
  reg [8:0] pointerOrCharacter_31; // @[treeGenerator.scala 29:31]
  reg [31:0] _RAND_63;
  reg  isCharacter_0; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_64;
  reg  isCharacter_1; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_65;
  reg  isCharacter_2; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_66;
  reg  isCharacter_3; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_67;
  reg  isCharacter_4; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_68;
  reg  isCharacter_5; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_69;
  reg  isCharacter_6; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_70;
  reg  isCharacter_7; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_71;
  reg  isCharacter_8; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_72;
  reg  isCharacter_9; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_73;
  reg  isCharacter_10; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_74;
  reg  isCharacter_11; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_75;
  reg  isCharacter_12; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_76;
  reg  isCharacter_13; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_77;
  reg  isCharacter_14; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_78;
  reg  isCharacter_15; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_79;
  reg  isCharacter_16; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_80;
  reg  isCharacter_17; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_81;
  reg  isCharacter_18; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_82;
  reg  isCharacter_19; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_83;
  reg  isCharacter_20; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_84;
  reg  isCharacter_21; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_85;
  reg  isCharacter_22; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_86;
  reg  isCharacter_23; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_87;
  reg  isCharacter_24; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_88;
  reg  isCharacter_25; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_89;
  reg  isCharacter_26; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_90;
  reg  isCharacter_27; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_91;
  reg  isCharacter_28; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_92;
  reg  isCharacter_29; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_93;
  reg  isCharacter_30; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_94;
  reg  isCharacter_31; // @[treeGenerator.scala 39:24]
  reg [31:0] _RAND_95;
  reg [12:0] newFrequency; // @[treeGenerator.scala 43:25]
  reg [31:0] _RAND_96;
  reg [8:0] newPointer; // @[treeGenerator.scala 44:23]
  reg [31:0] _RAND_97;
  reg [5:0] validRoots; // @[treeGenerator.scala 48:23]
  reg [31:0] _RAND_98;
  reg [8:0] leftNode_0; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_99;
  reg [8:0] leftNode_1; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_100;
  reg [8:0] leftNode_2; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_101;
  reg [8:0] leftNode_3; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_102;
  reg [8:0] leftNode_4; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_103;
  reg [8:0] leftNode_5; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_104;
  reg [8:0] leftNode_6; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_105;
  reg [8:0] leftNode_7; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_106;
  reg [8:0] leftNode_8; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_107;
  reg [8:0] leftNode_9; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_108;
  reg [8:0] leftNode_10; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_109;
  reg [8:0] leftNode_11; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_110;
  reg [8:0] leftNode_12; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_111;
  reg [8:0] leftNode_13; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_112;
  reg [8:0] leftNode_14; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_113;
  reg [8:0] leftNode_15; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_114;
  reg [8:0] leftNode_16; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_115;
  reg [8:0] leftNode_17; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_116;
  reg [8:0] leftNode_18; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_117;
  reg [8:0] leftNode_19; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_118;
  reg [8:0] leftNode_20; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_119;
  reg [8:0] leftNode_21; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_120;
  reg [8:0] leftNode_22; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_121;
  reg [8:0] leftNode_23; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_122;
  reg [8:0] leftNode_24; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_123;
  reg [8:0] leftNode_25; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_124;
  reg [8:0] leftNode_26; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_125;
  reg [8:0] leftNode_27; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_126;
  reg [8:0] leftNode_28; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_127;
  reg [8:0] leftNode_29; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_128;
  reg [8:0] leftNode_30; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_129;
  reg [8:0] leftNode_31; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_130;
  reg [8:0] leftNode_32; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_131;
  reg [8:0] leftNode_33; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_132;
  reg [8:0] leftNode_34; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_133;
  reg [8:0] leftNode_35; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_134;
  reg [8:0] leftNode_36; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_135;
  reg [8:0] leftNode_37; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_136;
  reg [8:0] leftNode_38; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_137;
  reg [8:0] leftNode_39; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_138;
  reg [8:0] leftNode_40; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_139;
  reg [8:0] leftNode_41; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_140;
  reg [8:0] leftNode_42; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_141;
  reg [8:0] leftNode_43; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_142;
  reg [8:0] leftNode_44; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_143;
  reg [8:0] leftNode_45; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_144;
  reg [8:0] leftNode_46; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_145;
  reg [8:0] leftNode_47; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_146;
  reg [8:0] leftNode_48; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_147;
  reg [8:0] leftNode_49; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_148;
  reg [8:0] leftNode_50; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_149;
  reg [8:0] leftNode_51; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_150;
  reg [8:0] leftNode_52; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_151;
  reg [8:0] leftNode_53; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_152;
  reg [8:0] leftNode_54; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_153;
  reg [8:0] leftNode_55; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_154;
  reg [8:0] leftNode_56; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_155;
  reg [8:0] leftNode_57; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_156;
  reg [8:0] leftNode_58; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_157;
  reg [8:0] leftNode_59; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_158;
  reg [8:0] leftNode_60; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_159;
  reg [8:0] leftNode_61; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_160;
  reg [8:0] leftNode_62; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_161;
  reg [8:0] leftNode_63; // @[treeGenerator.scala 54:21]
  reg [31:0] _RAND_162;
  reg [8:0] rightNode_0; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_163;
  reg [8:0] rightNode_1; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_164;
  reg [8:0] rightNode_2; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_165;
  reg [8:0] rightNode_3; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_166;
  reg [8:0] rightNode_4; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_167;
  reg [8:0] rightNode_5; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_168;
  reg [8:0] rightNode_6; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_169;
  reg [8:0] rightNode_7; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_170;
  reg [8:0] rightNode_8; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_171;
  reg [8:0] rightNode_9; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_172;
  reg [8:0] rightNode_10; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_173;
  reg [8:0] rightNode_11; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_174;
  reg [8:0] rightNode_12; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_175;
  reg [8:0] rightNode_13; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_176;
  reg [8:0] rightNode_14; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_177;
  reg [8:0] rightNode_15; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_178;
  reg [8:0] rightNode_16; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_179;
  reg [8:0] rightNode_17; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_180;
  reg [8:0] rightNode_18; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_181;
  reg [8:0] rightNode_19; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_182;
  reg [8:0] rightNode_20; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_183;
  reg [8:0] rightNode_21; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_184;
  reg [8:0] rightNode_22; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_185;
  reg [8:0] rightNode_23; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_186;
  reg [8:0] rightNode_24; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_187;
  reg [8:0] rightNode_25; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_188;
  reg [8:0] rightNode_26; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_189;
  reg [8:0] rightNode_27; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_190;
  reg [8:0] rightNode_28; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_191;
  reg [8:0] rightNode_29; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_192;
  reg [8:0] rightNode_30; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_193;
  reg [8:0] rightNode_31; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_194;
  reg [8:0] rightNode_32; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_195;
  reg [8:0] rightNode_33; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_196;
  reg [8:0] rightNode_34; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_197;
  reg [8:0] rightNode_35; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_198;
  reg [8:0] rightNode_36; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_199;
  reg [8:0] rightNode_37; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_200;
  reg [8:0] rightNode_38; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_201;
  reg [8:0] rightNode_39; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_202;
  reg [8:0] rightNode_40; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_203;
  reg [8:0] rightNode_41; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_204;
  reg [8:0] rightNode_42; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_205;
  reg [8:0] rightNode_43; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_206;
  reg [8:0] rightNode_44; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_207;
  reg [8:0] rightNode_45; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_208;
  reg [8:0] rightNode_46; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_209;
  reg [8:0] rightNode_47; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_210;
  reg [8:0] rightNode_48; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_211;
  reg [8:0] rightNode_49; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_212;
  reg [8:0] rightNode_50; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_213;
  reg [8:0] rightNode_51; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_214;
  reg [8:0] rightNode_52; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_215;
  reg [8:0] rightNode_53; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_216;
  reg [8:0] rightNode_54; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_217;
  reg [8:0] rightNode_55; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_218;
  reg [8:0] rightNode_56; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_219;
  reg [8:0] rightNode_57; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_220;
  reg [8:0] rightNode_58; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_221;
  reg [8:0] rightNode_59; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_222;
  reg [8:0] rightNode_60; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_223;
  reg [8:0] rightNode_61; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_224;
  reg [8:0] rightNode_62; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_225;
  reg [8:0] rightNode_63; // @[treeGenerator.scala 57:22]
  reg [31:0] _RAND_226;
  reg  leftNodeIsCharacter_0; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_227;
  reg  leftNodeIsCharacter_1; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_228;
  reg  leftNodeIsCharacter_2; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_229;
  reg  leftNodeIsCharacter_3; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_230;
  reg  leftNodeIsCharacter_4; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_231;
  reg  leftNodeIsCharacter_5; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_232;
  reg  leftNodeIsCharacter_6; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_233;
  reg  leftNodeIsCharacter_7; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_234;
  reg  leftNodeIsCharacter_8; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_235;
  reg  leftNodeIsCharacter_9; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_236;
  reg  leftNodeIsCharacter_10; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_237;
  reg  leftNodeIsCharacter_11; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_238;
  reg  leftNodeIsCharacter_12; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_239;
  reg  leftNodeIsCharacter_13; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_240;
  reg  leftNodeIsCharacter_14; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_241;
  reg  leftNodeIsCharacter_15; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_242;
  reg  leftNodeIsCharacter_16; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_243;
  reg  leftNodeIsCharacter_17; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_244;
  reg  leftNodeIsCharacter_18; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_245;
  reg  leftNodeIsCharacter_19; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_246;
  reg  leftNodeIsCharacter_20; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_247;
  reg  leftNodeIsCharacter_21; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_248;
  reg  leftNodeIsCharacter_22; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_249;
  reg  leftNodeIsCharacter_23; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_250;
  reg  leftNodeIsCharacter_24; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_251;
  reg  leftNodeIsCharacter_25; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_252;
  reg  leftNodeIsCharacter_26; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_253;
  reg  leftNodeIsCharacter_27; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_254;
  reg  leftNodeIsCharacter_28; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_255;
  reg  leftNodeIsCharacter_29; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_256;
  reg  leftNodeIsCharacter_30; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_257;
  reg  leftNodeIsCharacter_31; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_258;
  reg  leftNodeIsCharacter_32; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_259;
  reg  leftNodeIsCharacter_33; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_260;
  reg  leftNodeIsCharacter_34; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_261;
  reg  leftNodeIsCharacter_35; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_262;
  reg  leftNodeIsCharacter_36; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_263;
  reg  leftNodeIsCharacter_37; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_264;
  reg  leftNodeIsCharacter_38; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_265;
  reg  leftNodeIsCharacter_39; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_266;
  reg  leftNodeIsCharacter_40; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_267;
  reg  leftNodeIsCharacter_41; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_268;
  reg  leftNodeIsCharacter_42; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_269;
  reg  leftNodeIsCharacter_43; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_270;
  reg  leftNodeIsCharacter_44; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_271;
  reg  leftNodeIsCharacter_45; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_272;
  reg  leftNodeIsCharacter_46; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_273;
  reg  leftNodeIsCharacter_47; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_274;
  reg  leftNodeIsCharacter_48; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_275;
  reg  leftNodeIsCharacter_49; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_276;
  reg  leftNodeIsCharacter_50; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_277;
  reg  leftNodeIsCharacter_51; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_278;
  reg  leftNodeIsCharacter_52; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_279;
  reg  leftNodeIsCharacter_53; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_280;
  reg  leftNodeIsCharacter_54; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_281;
  reg  leftNodeIsCharacter_55; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_282;
  reg  leftNodeIsCharacter_56; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_283;
  reg  leftNodeIsCharacter_57; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_284;
  reg  leftNodeIsCharacter_58; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_285;
  reg  leftNodeIsCharacter_59; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_286;
  reg  leftNodeIsCharacter_60; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_287;
  reg  leftNodeIsCharacter_61; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_288;
  reg  leftNodeIsCharacter_62; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_289;
  reg  leftNodeIsCharacter_63; // @[treeGenerator.scala 60:32]
  reg [31:0] _RAND_290;
  reg  rightNodeIsCharacter_0; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_291;
  reg  rightNodeIsCharacter_1; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_292;
  reg  rightNodeIsCharacter_2; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_293;
  reg  rightNodeIsCharacter_3; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_294;
  reg  rightNodeIsCharacter_4; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_295;
  reg  rightNodeIsCharacter_5; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_296;
  reg  rightNodeIsCharacter_6; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_297;
  reg  rightNodeIsCharacter_7; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_298;
  reg  rightNodeIsCharacter_8; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_299;
  reg  rightNodeIsCharacter_9; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_300;
  reg  rightNodeIsCharacter_10; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_301;
  reg  rightNodeIsCharacter_11; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_302;
  reg  rightNodeIsCharacter_12; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_303;
  reg  rightNodeIsCharacter_13; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_304;
  reg  rightNodeIsCharacter_14; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_305;
  reg  rightNodeIsCharacter_15; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_306;
  reg  rightNodeIsCharacter_16; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_307;
  reg  rightNodeIsCharacter_17; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_308;
  reg  rightNodeIsCharacter_18; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_309;
  reg  rightNodeIsCharacter_19; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_310;
  reg  rightNodeIsCharacter_20; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_311;
  reg  rightNodeIsCharacter_21; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_312;
  reg  rightNodeIsCharacter_22; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_313;
  reg  rightNodeIsCharacter_23; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_314;
  reg  rightNodeIsCharacter_24; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_315;
  reg  rightNodeIsCharacter_25; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_316;
  reg  rightNodeIsCharacter_26; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_317;
  reg  rightNodeIsCharacter_27; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_318;
  reg  rightNodeIsCharacter_28; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_319;
  reg  rightNodeIsCharacter_29; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_320;
  reg  rightNodeIsCharacter_30; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_321;
  reg  rightNodeIsCharacter_31; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_322;
  reg  rightNodeIsCharacter_32; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_323;
  reg  rightNodeIsCharacter_33; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_324;
  reg  rightNodeIsCharacter_34; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_325;
  reg  rightNodeIsCharacter_35; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_326;
  reg  rightNodeIsCharacter_36; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_327;
  reg  rightNodeIsCharacter_37; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_328;
  reg  rightNodeIsCharacter_38; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_329;
  reg  rightNodeIsCharacter_39; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_330;
  reg  rightNodeIsCharacter_40; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_331;
  reg  rightNodeIsCharacter_41; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_332;
  reg  rightNodeIsCharacter_42; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_333;
  reg  rightNodeIsCharacter_43; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_334;
  reg  rightNodeIsCharacter_44; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_335;
  reg  rightNodeIsCharacter_45; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_336;
  reg  rightNodeIsCharacter_46; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_337;
  reg  rightNodeIsCharacter_47; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_338;
  reg  rightNodeIsCharacter_48; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_339;
  reg  rightNodeIsCharacter_49; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_340;
  reg  rightNodeIsCharacter_50; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_341;
  reg  rightNodeIsCharacter_51; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_342;
  reg  rightNodeIsCharacter_52; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_343;
  reg  rightNodeIsCharacter_53; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_344;
  reg  rightNodeIsCharacter_54; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_345;
  reg  rightNodeIsCharacter_55; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_346;
  reg  rightNodeIsCharacter_56; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_347;
  reg  rightNodeIsCharacter_57; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_348;
  reg  rightNodeIsCharacter_58; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_349;
  reg  rightNodeIsCharacter_59; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_350;
  reg  rightNodeIsCharacter_60; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_351;
  reg  rightNodeIsCharacter_61; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_352;
  reg  rightNodeIsCharacter_62; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_353;
  reg  rightNodeIsCharacter_63; // @[treeGenerator.scala 61:33]
  reg [31:0] _RAND_354;
  reg [5:0] upperNodeIndex; // @[treeGenerator.scala 65:27]
  reg [31:0] _RAND_355;
  reg [5:0] lowerNodeIndex; // @[treeGenerator.scala 66:27]
  reg [31:0] _RAND_356;
  reg [6:0] validNodes; // @[treeGenerator.scala 71:23]
  reg [31:0] _RAND_357;
  reg [5:0] validCharacters; // @[treeGenerator.scala 75:28]
  reg [31:0] _RAND_358;
  wire  nonZeroFrequencies_0 = io_inputs_sortedFrequency_0 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_1 = io_inputs_sortedFrequency_1 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_2 = io_inputs_sortedFrequency_2 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_3 = io_inputs_sortedFrequency_3 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_4 = io_inputs_sortedFrequency_4 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_5 = io_inputs_sortedFrequency_5 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_6 = io_inputs_sortedFrequency_6 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_7 = io_inputs_sortedFrequency_7 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_8 = io_inputs_sortedFrequency_8 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_9 = io_inputs_sortedFrequency_9 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_10 = io_inputs_sortedFrequency_10 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_11 = io_inputs_sortedFrequency_11 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_12 = io_inputs_sortedFrequency_12 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_13 = io_inputs_sortedFrequency_13 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_14 = io_inputs_sortedFrequency_14 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_15 = io_inputs_sortedFrequency_15 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_16 = io_inputs_sortedFrequency_16 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_17 = io_inputs_sortedFrequency_17 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_18 = io_inputs_sortedFrequency_18 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_19 = io_inputs_sortedFrequency_19 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_20 = io_inputs_sortedFrequency_20 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_21 = io_inputs_sortedFrequency_21 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_22 = io_inputs_sortedFrequency_22 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_23 = io_inputs_sortedFrequency_23 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_24 = io_inputs_sortedFrequency_24 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_25 = io_inputs_sortedFrequency_25 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_26 = io_inputs_sortedFrequency_26 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_27 = io_inputs_sortedFrequency_27 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_28 = io_inputs_sortedFrequency_28 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_29 = io_inputs_sortedFrequency_29 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_30 = io_inputs_sortedFrequency_30 != 13'h0; // @[treeGenerator.scala 81:67]
  wire  nonZeroFrequencies_31 = io_inputs_sortedFrequency_31 != 13'h0; // @[treeGenerator.scala 81:67]
  reg [1:0] state; // @[treeGenerator.scala 94:22]
  reg [31:0] _RAND_359;
  wire  _T_32 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire [7:0] _T_40 = {nonZeroFrequencies_7,nonZeroFrequencies_6,nonZeroFrequencies_5,nonZeroFrequencies_4,nonZeroFrequencies_3,nonZeroFrequencies_2,nonZeroFrequencies_1,nonZeroFrequencies_0}; // @[treeGenerator.scala 105:57]
  wire [15:0] _T_48 = {nonZeroFrequencies_15,nonZeroFrequencies_14,nonZeroFrequencies_13,nonZeroFrequencies_12,nonZeroFrequencies_11,nonZeroFrequencies_10,nonZeroFrequencies_9,nonZeroFrequencies_8,_T_40}; // @[treeGenerator.scala 105:57]
  wire [7:0] _T_55 = {nonZeroFrequencies_23,nonZeroFrequencies_22,nonZeroFrequencies_21,nonZeroFrequencies_20,nonZeroFrequencies_19,nonZeroFrequencies_18,nonZeroFrequencies_17,nonZeroFrequencies_16}; // @[treeGenerator.scala 105:57]
  wire [31:0] _T_64 = {nonZeroFrequencies_31,nonZeroFrequencies_30,nonZeroFrequencies_29,nonZeroFrequencies_28,nonZeroFrequencies_27,nonZeroFrequencies_26,nonZeroFrequencies_25,nonZeroFrequencies_24,_T_55,_T_48}; // @[treeGenerator.scala 105:57]
  wire [1:0] _T_97 = _T_64[0] + _T_64[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_99 = _T_64[2] + _T_64[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_101 = _T_97 + _T_99; // @[Bitwise.scala 47:55]
  wire [1:0] _T_103 = _T_64[4] + _T_64[5]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_105 = _T_64[6] + _T_64[7]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_107 = _T_103 + _T_105; // @[Bitwise.scala 47:55]
  wire [3:0] _T_109 = _T_101 + _T_107; // @[Bitwise.scala 47:55]
  wire [1:0] _T_111 = _T_64[8] + _T_64[9]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_113 = _T_64[10] + _T_64[11]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_115 = _T_111 + _T_113; // @[Bitwise.scala 47:55]
  wire [1:0] _T_117 = _T_64[12] + _T_64[13]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_119 = _T_64[14] + _T_64[15]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_121 = _T_117 + _T_119; // @[Bitwise.scala 47:55]
  wire [3:0] _T_123 = _T_115 + _T_121; // @[Bitwise.scala 47:55]
  wire [4:0] _T_125 = _T_109 + _T_123; // @[Bitwise.scala 47:55]
  wire [1:0] _T_127 = _T_64[16] + _T_64[17]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_129 = _T_64[18] + _T_64[19]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_131 = _T_127 + _T_129; // @[Bitwise.scala 47:55]
  wire [1:0] _T_133 = _T_64[20] + _T_64[21]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_135 = _T_64[22] + _T_64[23]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_137 = _T_133 + _T_135; // @[Bitwise.scala 47:55]
  wire [3:0] _T_139 = _T_131 + _T_137; // @[Bitwise.scala 47:55]
  wire [1:0] _T_141 = _T_64[24] + _T_64[25]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_143 = _T_64[26] + _T_64[27]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_145 = _T_141 + _T_143; // @[Bitwise.scala 47:55]
  wire [1:0] _T_147 = _T_64[28] + _T_64[29]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_149 = _T_64[30] + _T_64[31]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_151 = _T_147 + _T_149; // @[Bitwise.scala 47:55]
  wire [3:0] _T_153 = _T_145 + _T_151; // @[Bitwise.scala 47:55]
  wire [4:0] _T_155 = _T_139 + _T_153; // @[Bitwise.scala 47:55]
  wire [5:0] _T_157 = _T_125 + _T_155; // @[Bitwise.scala 47:55]
  wire  _GEN_66 = io_start | isCharacter_0; // @[treeGenerator.scala 98:22]
  wire  _GEN_67 = io_start | isCharacter_1; // @[treeGenerator.scala 98:22]
  wire  _GEN_68 = io_start | isCharacter_2; // @[treeGenerator.scala 98:22]
  wire  _GEN_69 = io_start | isCharacter_3; // @[treeGenerator.scala 98:22]
  wire  _GEN_70 = io_start | isCharacter_4; // @[treeGenerator.scala 98:22]
  wire  _GEN_71 = io_start | isCharacter_5; // @[treeGenerator.scala 98:22]
  wire  _GEN_72 = io_start | isCharacter_6; // @[treeGenerator.scala 98:22]
  wire  _GEN_73 = io_start | isCharacter_7; // @[treeGenerator.scala 98:22]
  wire  _GEN_74 = io_start | isCharacter_8; // @[treeGenerator.scala 98:22]
  wire  _GEN_75 = io_start | isCharacter_9; // @[treeGenerator.scala 98:22]
  wire  _GEN_76 = io_start | isCharacter_10; // @[treeGenerator.scala 98:22]
  wire  _GEN_77 = io_start | isCharacter_11; // @[treeGenerator.scala 98:22]
  wire  _GEN_78 = io_start | isCharacter_12; // @[treeGenerator.scala 98:22]
  wire  _GEN_79 = io_start | isCharacter_13; // @[treeGenerator.scala 98:22]
  wire  _GEN_80 = io_start | isCharacter_14; // @[treeGenerator.scala 98:22]
  wire  _GEN_81 = io_start | isCharacter_15; // @[treeGenerator.scala 98:22]
  wire  _GEN_82 = io_start | isCharacter_16; // @[treeGenerator.scala 98:22]
  wire  _GEN_83 = io_start | isCharacter_17; // @[treeGenerator.scala 98:22]
  wire  _GEN_84 = io_start | isCharacter_18; // @[treeGenerator.scala 98:22]
  wire  _GEN_85 = io_start | isCharacter_19; // @[treeGenerator.scala 98:22]
  wire  _GEN_86 = io_start | isCharacter_20; // @[treeGenerator.scala 98:22]
  wire  _GEN_87 = io_start | isCharacter_21; // @[treeGenerator.scala 98:22]
  wire  _GEN_88 = io_start | isCharacter_22; // @[treeGenerator.scala 98:22]
  wire  _GEN_89 = io_start | isCharacter_23; // @[treeGenerator.scala 98:22]
  wire  _GEN_90 = io_start | isCharacter_24; // @[treeGenerator.scala 98:22]
  wire  _GEN_91 = io_start | isCharacter_25; // @[treeGenerator.scala 98:22]
  wire  _GEN_92 = io_start | isCharacter_26; // @[treeGenerator.scala 98:22]
  wire  _GEN_93 = io_start | isCharacter_27; // @[treeGenerator.scala 98:22]
  wire  _GEN_94 = io_start | isCharacter_28; // @[treeGenerator.scala 98:22]
  wire  _GEN_95 = io_start | isCharacter_29; // @[treeGenerator.scala 98:22]
  wire  _GEN_96 = io_start | isCharacter_30; // @[treeGenerator.scala 98:22]
  wire  _GEN_97 = io_start | isCharacter_31; // @[treeGenerator.scala 98:22]
  wire  _T_284 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_285 = validRoots < 6'h2; // @[treeGenerator.scala 111:23]
  wire  _T_286 = validNodes == 7'h0; // @[treeGenerator.scala 112:25]
  wire  _GEN_103 = _T_286 | leftNodeIsCharacter_0; // @[treeGenerator.scala 112:34]
  wire [6:0] _T_288 = validNodes + 7'h1; // @[treeGenerator.scala 128:34]
  wire [5:0] _T_290 = validRoots - 6'h1; // @[treeGenerator.scala 129:34]
  wire [5:0] _T_293 = validRoots - 6'h2; // @[treeGenerator.scala 130:63]
  wire [8:0] _GEN_169 = 5'h1 == _T_293[4:0] ? pointerOrCharacter_1 : pointerOrCharacter_0; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_170 = 5'h2 == _T_293[4:0] ? pointerOrCharacter_2 : _GEN_169; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_171 = 5'h3 == _T_293[4:0] ? pointerOrCharacter_3 : _GEN_170; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_172 = 5'h4 == _T_293[4:0] ? pointerOrCharacter_4 : _GEN_171; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_173 = 5'h5 == _T_293[4:0] ? pointerOrCharacter_5 : _GEN_172; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_174 = 5'h6 == _T_293[4:0] ? pointerOrCharacter_6 : _GEN_173; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_175 = 5'h7 == _T_293[4:0] ? pointerOrCharacter_7 : _GEN_174; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_176 = 5'h8 == _T_293[4:0] ? pointerOrCharacter_8 : _GEN_175; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_177 = 5'h9 == _T_293[4:0] ? pointerOrCharacter_9 : _GEN_176; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_178 = 5'ha == _T_293[4:0] ? pointerOrCharacter_10 : _GEN_177; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_179 = 5'hb == _T_293[4:0] ? pointerOrCharacter_11 : _GEN_178; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_180 = 5'hc == _T_293[4:0] ? pointerOrCharacter_12 : _GEN_179; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_181 = 5'hd == _T_293[4:0] ? pointerOrCharacter_13 : _GEN_180; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_182 = 5'he == _T_293[4:0] ? pointerOrCharacter_14 : _GEN_181; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_183 = 5'hf == _T_293[4:0] ? pointerOrCharacter_15 : _GEN_182; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_184 = 5'h10 == _T_293[4:0] ? pointerOrCharacter_16 : _GEN_183; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_185 = 5'h11 == _T_293[4:0] ? pointerOrCharacter_17 : _GEN_184; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_186 = 5'h12 == _T_293[4:0] ? pointerOrCharacter_18 : _GEN_185; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_187 = 5'h13 == _T_293[4:0] ? pointerOrCharacter_19 : _GEN_186; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_188 = 5'h14 == _T_293[4:0] ? pointerOrCharacter_20 : _GEN_187; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_189 = 5'h15 == _T_293[4:0] ? pointerOrCharacter_21 : _GEN_188; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_190 = 5'h16 == _T_293[4:0] ? pointerOrCharacter_22 : _GEN_189; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_191 = 5'h17 == _T_293[4:0] ? pointerOrCharacter_23 : _GEN_190; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_192 = 5'h18 == _T_293[4:0] ? pointerOrCharacter_24 : _GEN_191; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_193 = 5'h19 == _T_293[4:0] ? pointerOrCharacter_25 : _GEN_192; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_194 = 5'h1a == _T_293[4:0] ? pointerOrCharacter_26 : _GEN_193; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_195 = 5'h1b == _T_293[4:0] ? pointerOrCharacter_27 : _GEN_194; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_196 = 5'h1c == _T_293[4:0] ? pointerOrCharacter_28 : _GEN_195; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_197 = 5'h1d == _T_293[4:0] ? pointerOrCharacter_29 : _GEN_196; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_198 = 5'h1e == _T_293[4:0] ? pointerOrCharacter_30 : _GEN_197; // @[treeGenerator.scala 130:30]
  wire [8:0] _GEN_199 = 5'h1f == _T_293[4:0] ? pointerOrCharacter_31 : _GEN_198; // @[treeGenerator.scala 130:30]
  wire  _GEN_265 = 5'h1 == _T_293[4:0] ? isCharacter_1 : isCharacter_0; // @[treeGenerator.scala 131:41]
  wire  _GEN_266 = 5'h2 == _T_293[4:0] ? isCharacter_2 : _GEN_265; // @[treeGenerator.scala 131:41]
  wire  _GEN_267 = 5'h3 == _T_293[4:0] ? isCharacter_3 : _GEN_266; // @[treeGenerator.scala 131:41]
  wire  _GEN_268 = 5'h4 == _T_293[4:0] ? isCharacter_4 : _GEN_267; // @[treeGenerator.scala 131:41]
  wire  _GEN_269 = 5'h5 == _T_293[4:0] ? isCharacter_5 : _GEN_268; // @[treeGenerator.scala 131:41]
  wire  _GEN_270 = 5'h6 == _T_293[4:0] ? isCharacter_6 : _GEN_269; // @[treeGenerator.scala 131:41]
  wire  _GEN_271 = 5'h7 == _T_293[4:0] ? isCharacter_7 : _GEN_270; // @[treeGenerator.scala 131:41]
  wire  _GEN_272 = 5'h8 == _T_293[4:0] ? isCharacter_8 : _GEN_271; // @[treeGenerator.scala 131:41]
  wire  _GEN_273 = 5'h9 == _T_293[4:0] ? isCharacter_9 : _GEN_272; // @[treeGenerator.scala 131:41]
  wire  _GEN_274 = 5'ha == _T_293[4:0] ? isCharacter_10 : _GEN_273; // @[treeGenerator.scala 131:41]
  wire  _GEN_275 = 5'hb == _T_293[4:0] ? isCharacter_11 : _GEN_274; // @[treeGenerator.scala 131:41]
  wire  _GEN_276 = 5'hc == _T_293[4:0] ? isCharacter_12 : _GEN_275; // @[treeGenerator.scala 131:41]
  wire  _GEN_277 = 5'hd == _T_293[4:0] ? isCharacter_13 : _GEN_276; // @[treeGenerator.scala 131:41]
  wire  _GEN_278 = 5'he == _T_293[4:0] ? isCharacter_14 : _GEN_277; // @[treeGenerator.scala 131:41]
  wire  _GEN_279 = 5'hf == _T_293[4:0] ? isCharacter_15 : _GEN_278; // @[treeGenerator.scala 131:41]
  wire  _GEN_280 = 5'h10 == _T_293[4:0] ? isCharacter_16 : _GEN_279; // @[treeGenerator.scala 131:41]
  wire  _GEN_281 = 5'h11 == _T_293[4:0] ? isCharacter_17 : _GEN_280; // @[treeGenerator.scala 131:41]
  wire  _GEN_282 = 5'h12 == _T_293[4:0] ? isCharacter_18 : _GEN_281; // @[treeGenerator.scala 131:41]
  wire  _GEN_283 = 5'h13 == _T_293[4:0] ? isCharacter_19 : _GEN_282; // @[treeGenerator.scala 131:41]
  wire  _GEN_284 = 5'h14 == _T_293[4:0] ? isCharacter_20 : _GEN_283; // @[treeGenerator.scala 131:41]
  wire  _GEN_285 = 5'h15 == _T_293[4:0] ? isCharacter_21 : _GEN_284; // @[treeGenerator.scala 131:41]
  wire  _GEN_286 = 5'h16 == _T_293[4:0] ? isCharacter_22 : _GEN_285; // @[treeGenerator.scala 131:41]
  wire  _GEN_287 = 5'h17 == _T_293[4:0] ? isCharacter_23 : _GEN_286; // @[treeGenerator.scala 131:41]
  wire  _GEN_288 = 5'h18 == _T_293[4:0] ? isCharacter_24 : _GEN_287; // @[treeGenerator.scala 131:41]
  wire  _GEN_289 = 5'h19 == _T_293[4:0] ? isCharacter_25 : _GEN_288; // @[treeGenerator.scala 131:41]
  wire  _GEN_290 = 5'h1a == _T_293[4:0] ? isCharacter_26 : _GEN_289; // @[treeGenerator.scala 131:41]
  wire  _GEN_291 = 5'h1b == _T_293[4:0] ? isCharacter_27 : _GEN_290; // @[treeGenerator.scala 131:41]
  wire  _GEN_292 = 5'h1c == _T_293[4:0] ? isCharacter_28 : _GEN_291; // @[treeGenerator.scala 131:41]
  wire  _GEN_293 = 5'h1d == _T_293[4:0] ? isCharacter_29 : _GEN_292; // @[treeGenerator.scala 131:41]
  wire  _GEN_294 = 5'h1e == _T_293[4:0] ? isCharacter_30 : _GEN_293; // @[treeGenerator.scala 131:41]
  wire  _GEN_295 = 5'h1f == _T_293[4:0] ? isCharacter_31 : _GEN_294; // @[treeGenerator.scala 131:41]
  wire [8:0] _GEN_361 = 5'h1 == _T_290[4:0] ? pointerOrCharacter_1 : pointerOrCharacter_0; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_362 = 5'h2 == _T_290[4:0] ? pointerOrCharacter_2 : _GEN_361; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_363 = 5'h3 == _T_290[4:0] ? pointerOrCharacter_3 : _GEN_362; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_364 = 5'h4 == _T_290[4:0] ? pointerOrCharacter_4 : _GEN_363; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_365 = 5'h5 == _T_290[4:0] ? pointerOrCharacter_5 : _GEN_364; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_366 = 5'h6 == _T_290[4:0] ? pointerOrCharacter_6 : _GEN_365; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_367 = 5'h7 == _T_290[4:0] ? pointerOrCharacter_7 : _GEN_366; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_368 = 5'h8 == _T_290[4:0] ? pointerOrCharacter_8 : _GEN_367; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_369 = 5'h9 == _T_290[4:0] ? pointerOrCharacter_9 : _GEN_368; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_370 = 5'ha == _T_290[4:0] ? pointerOrCharacter_10 : _GEN_369; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_371 = 5'hb == _T_290[4:0] ? pointerOrCharacter_11 : _GEN_370; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_372 = 5'hc == _T_290[4:0] ? pointerOrCharacter_12 : _GEN_371; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_373 = 5'hd == _T_290[4:0] ? pointerOrCharacter_13 : _GEN_372; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_374 = 5'he == _T_290[4:0] ? pointerOrCharacter_14 : _GEN_373; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_375 = 5'hf == _T_290[4:0] ? pointerOrCharacter_15 : _GEN_374; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_376 = 5'h10 == _T_290[4:0] ? pointerOrCharacter_16 : _GEN_375; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_377 = 5'h11 == _T_290[4:0] ? pointerOrCharacter_17 : _GEN_376; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_378 = 5'h12 == _T_290[4:0] ? pointerOrCharacter_18 : _GEN_377; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_379 = 5'h13 == _T_290[4:0] ? pointerOrCharacter_19 : _GEN_378; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_380 = 5'h14 == _T_290[4:0] ? pointerOrCharacter_20 : _GEN_379; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_381 = 5'h15 == _T_290[4:0] ? pointerOrCharacter_21 : _GEN_380; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_382 = 5'h16 == _T_290[4:0] ? pointerOrCharacter_22 : _GEN_381; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_383 = 5'h17 == _T_290[4:0] ? pointerOrCharacter_23 : _GEN_382; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_384 = 5'h18 == _T_290[4:0] ? pointerOrCharacter_24 : _GEN_383; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_385 = 5'h19 == _T_290[4:0] ? pointerOrCharacter_25 : _GEN_384; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_386 = 5'h1a == _T_290[4:0] ? pointerOrCharacter_26 : _GEN_385; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_387 = 5'h1b == _T_290[4:0] ? pointerOrCharacter_27 : _GEN_386; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_388 = 5'h1c == _T_290[4:0] ? pointerOrCharacter_28 : _GEN_387; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_389 = 5'h1d == _T_290[4:0] ? pointerOrCharacter_29 : _GEN_388; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_390 = 5'h1e == _T_290[4:0] ? pointerOrCharacter_30 : _GEN_389; // @[treeGenerator.scala 132:31]
  wire [8:0] _GEN_391 = 5'h1f == _T_290[4:0] ? pointerOrCharacter_31 : _GEN_390; // @[treeGenerator.scala 132:31]
  wire  _GEN_457 = 5'h1 == _T_290[4:0] ? isCharacter_1 : isCharacter_0; // @[treeGenerator.scala 133:42]
  wire  _GEN_458 = 5'h2 == _T_290[4:0] ? isCharacter_2 : _GEN_457; // @[treeGenerator.scala 133:42]
  wire  _GEN_459 = 5'h3 == _T_290[4:0] ? isCharacter_3 : _GEN_458; // @[treeGenerator.scala 133:42]
  wire  _GEN_460 = 5'h4 == _T_290[4:0] ? isCharacter_4 : _GEN_459; // @[treeGenerator.scala 133:42]
  wire  _GEN_461 = 5'h5 == _T_290[4:0] ? isCharacter_5 : _GEN_460; // @[treeGenerator.scala 133:42]
  wire  _GEN_462 = 5'h6 == _T_290[4:0] ? isCharacter_6 : _GEN_461; // @[treeGenerator.scala 133:42]
  wire  _GEN_463 = 5'h7 == _T_290[4:0] ? isCharacter_7 : _GEN_462; // @[treeGenerator.scala 133:42]
  wire  _GEN_464 = 5'h8 == _T_290[4:0] ? isCharacter_8 : _GEN_463; // @[treeGenerator.scala 133:42]
  wire  _GEN_465 = 5'h9 == _T_290[4:0] ? isCharacter_9 : _GEN_464; // @[treeGenerator.scala 133:42]
  wire  _GEN_466 = 5'ha == _T_290[4:0] ? isCharacter_10 : _GEN_465; // @[treeGenerator.scala 133:42]
  wire  _GEN_467 = 5'hb == _T_290[4:0] ? isCharacter_11 : _GEN_466; // @[treeGenerator.scala 133:42]
  wire  _GEN_468 = 5'hc == _T_290[4:0] ? isCharacter_12 : _GEN_467; // @[treeGenerator.scala 133:42]
  wire  _GEN_469 = 5'hd == _T_290[4:0] ? isCharacter_13 : _GEN_468; // @[treeGenerator.scala 133:42]
  wire  _GEN_470 = 5'he == _T_290[4:0] ? isCharacter_14 : _GEN_469; // @[treeGenerator.scala 133:42]
  wire  _GEN_471 = 5'hf == _T_290[4:0] ? isCharacter_15 : _GEN_470; // @[treeGenerator.scala 133:42]
  wire  _GEN_472 = 5'h10 == _T_290[4:0] ? isCharacter_16 : _GEN_471; // @[treeGenerator.scala 133:42]
  wire  _GEN_473 = 5'h11 == _T_290[4:0] ? isCharacter_17 : _GEN_472; // @[treeGenerator.scala 133:42]
  wire  _GEN_474 = 5'h12 == _T_290[4:0] ? isCharacter_18 : _GEN_473; // @[treeGenerator.scala 133:42]
  wire  _GEN_475 = 5'h13 == _T_290[4:0] ? isCharacter_19 : _GEN_474; // @[treeGenerator.scala 133:42]
  wire  _GEN_476 = 5'h14 == _T_290[4:0] ? isCharacter_20 : _GEN_475; // @[treeGenerator.scala 133:42]
  wire  _GEN_477 = 5'h15 == _T_290[4:0] ? isCharacter_21 : _GEN_476; // @[treeGenerator.scala 133:42]
  wire  _GEN_478 = 5'h16 == _T_290[4:0] ? isCharacter_22 : _GEN_477; // @[treeGenerator.scala 133:42]
  wire  _GEN_479 = 5'h17 == _T_290[4:0] ? isCharacter_23 : _GEN_478; // @[treeGenerator.scala 133:42]
  wire  _GEN_480 = 5'h18 == _T_290[4:0] ? isCharacter_24 : _GEN_479; // @[treeGenerator.scala 133:42]
  wire  _GEN_481 = 5'h19 == _T_290[4:0] ? isCharacter_25 : _GEN_480; // @[treeGenerator.scala 133:42]
  wire  _GEN_482 = 5'h1a == _T_290[4:0] ? isCharacter_26 : _GEN_481; // @[treeGenerator.scala 133:42]
  wire  _GEN_483 = 5'h1b == _T_290[4:0] ? isCharacter_27 : _GEN_482; // @[treeGenerator.scala 133:42]
  wire  _GEN_484 = 5'h1c == _T_290[4:0] ? isCharacter_28 : _GEN_483; // @[treeGenerator.scala 133:42]
  wire  _GEN_485 = 5'h1d == _T_290[4:0] ? isCharacter_29 : _GEN_484; // @[treeGenerator.scala 133:42]
  wire  _GEN_486 = 5'h1e == _T_290[4:0] ? isCharacter_30 : _GEN_485; // @[treeGenerator.scala 133:42]
  wire  _GEN_487 = 5'h1f == _T_290[4:0] ? isCharacter_31 : _GEN_486; // @[treeGenerator.scala 133:42]
  wire [12:0] _GEN_489 = 5'h1 == _T_293[4:0] ? frequency_1 : frequency_0; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_490 = 5'h2 == _T_293[4:0] ? frequency_2 : _GEN_489; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_491 = 5'h3 == _T_293[4:0] ? frequency_3 : _GEN_490; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_492 = 5'h4 == _T_293[4:0] ? frequency_4 : _GEN_491; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_493 = 5'h5 == _T_293[4:0] ? frequency_5 : _GEN_492; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_494 = 5'h6 == _T_293[4:0] ? frequency_6 : _GEN_493; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_495 = 5'h7 == _T_293[4:0] ? frequency_7 : _GEN_494; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_496 = 5'h8 == _T_293[4:0] ? frequency_8 : _GEN_495; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_497 = 5'h9 == _T_293[4:0] ? frequency_9 : _GEN_496; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_498 = 5'ha == _T_293[4:0] ? frequency_10 : _GEN_497; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_499 = 5'hb == _T_293[4:0] ? frequency_11 : _GEN_498; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_500 = 5'hc == _T_293[4:0] ? frequency_12 : _GEN_499; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_501 = 5'hd == _T_293[4:0] ? frequency_13 : _GEN_500; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_502 = 5'he == _T_293[4:0] ? frequency_14 : _GEN_501; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_503 = 5'hf == _T_293[4:0] ? frequency_15 : _GEN_502; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_504 = 5'h10 == _T_293[4:0] ? frequency_16 : _GEN_503; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_505 = 5'h11 == _T_293[4:0] ? frequency_17 : _GEN_504; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_506 = 5'h12 == _T_293[4:0] ? frequency_18 : _GEN_505; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_507 = 5'h13 == _T_293[4:0] ? frequency_19 : _GEN_506; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_508 = 5'h14 == _T_293[4:0] ? frequency_20 : _GEN_507; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_509 = 5'h15 == _T_293[4:0] ? frequency_21 : _GEN_508; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_510 = 5'h16 == _T_293[4:0] ? frequency_22 : _GEN_509; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_511 = 5'h17 == _T_293[4:0] ? frequency_23 : _GEN_510; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_512 = 5'h18 == _T_293[4:0] ? frequency_24 : _GEN_511; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_513 = 5'h19 == _T_293[4:0] ? frequency_25 : _GEN_512; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_514 = 5'h1a == _T_293[4:0] ? frequency_26 : _GEN_513; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_515 = 5'h1b == _T_293[4:0] ? frequency_27 : _GEN_514; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_516 = 5'h1c == _T_293[4:0] ? frequency_28 : _GEN_515; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_517 = 5'h1d == _T_293[4:0] ? frequency_29 : _GEN_516; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_518 = 5'h1e == _T_293[4:0] ? frequency_30 : _GEN_517; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_519 = 5'h1f == _T_293[4:0] ? frequency_31 : _GEN_518; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_521 = 5'h1 == _T_290[4:0] ? frequency_1 : frequency_0; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_522 = 5'h2 == _T_290[4:0] ? frequency_2 : _GEN_521; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_523 = 5'h3 == _T_290[4:0] ? frequency_3 : _GEN_522; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_524 = 5'h4 == _T_290[4:0] ? frequency_4 : _GEN_523; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_525 = 5'h5 == _T_290[4:0] ? frequency_5 : _GEN_524; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_526 = 5'h6 == _T_290[4:0] ? frequency_6 : _GEN_525; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_527 = 5'h7 == _T_290[4:0] ? frequency_7 : _GEN_526; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_528 = 5'h8 == _T_290[4:0] ? frequency_8 : _GEN_527; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_529 = 5'h9 == _T_290[4:0] ? frequency_9 : _GEN_528; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_530 = 5'ha == _T_290[4:0] ? frequency_10 : _GEN_529; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_531 = 5'hb == _T_290[4:0] ? frequency_11 : _GEN_530; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_532 = 5'hc == _T_290[4:0] ? frequency_12 : _GEN_531; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_533 = 5'hd == _T_290[4:0] ? frequency_13 : _GEN_532; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_534 = 5'he == _T_290[4:0] ? frequency_14 : _GEN_533; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_535 = 5'hf == _T_290[4:0] ? frequency_15 : _GEN_534; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_536 = 5'h10 == _T_290[4:0] ? frequency_16 : _GEN_535; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_537 = 5'h11 == _T_290[4:0] ? frequency_17 : _GEN_536; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_538 = 5'h12 == _T_290[4:0] ? frequency_18 : _GEN_537; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_539 = 5'h13 == _T_290[4:0] ? frequency_19 : _GEN_538; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_540 = 5'h14 == _T_290[4:0] ? frequency_20 : _GEN_539; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_541 = 5'h15 == _T_290[4:0] ? frequency_21 : _GEN_540; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_542 = 5'h16 == _T_290[4:0] ? frequency_22 : _GEN_541; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_543 = 5'h17 == _T_290[4:0] ? frequency_23 : _GEN_542; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_544 = 5'h18 == _T_290[4:0] ? frequency_24 : _GEN_543; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_545 = 5'h19 == _T_290[4:0] ? frequency_25 : _GEN_544; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_546 = 5'h1a == _T_290[4:0] ? frequency_26 : _GEN_545; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_547 = 5'h1b == _T_290[4:0] ? frequency_27 : _GEN_546; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_548 = 5'h1c == _T_290[4:0] ? frequency_28 : _GEN_547; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_549 = 5'h1d == _T_290[4:0] ? frequency_29 : _GEN_548; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_550 = 5'h1e == _T_290[4:0] ? frequency_30 : _GEN_549; // @[treeGenerator.scala 140:53]
  wire [12:0] _GEN_551 = 5'h1f == _T_290[4:0] ? frequency_31 : _GEN_550; // @[treeGenerator.scala 140:53]
  wire [12:0] _T_314 = _GEN_519 + _GEN_551; // @[treeGenerator.scala 140:53]
  wire  _T_317 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_318 = upperNodeIndex == lowerNodeIndex; // @[treeGenerator.scala 152:25]
  wire [12:0] _GEN_817 = 5'h1 == upperNodeIndex[4:0] ? frequency_1 : frequency_0; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_818 = 5'h2 == upperNodeIndex[4:0] ? frequency_2 : _GEN_817; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_819 = 5'h3 == upperNodeIndex[4:0] ? frequency_3 : _GEN_818; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_820 = 5'h4 == upperNodeIndex[4:0] ? frequency_4 : _GEN_819; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_821 = 5'h5 == upperNodeIndex[4:0] ? frequency_5 : _GEN_820; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_822 = 5'h6 == upperNodeIndex[4:0] ? frequency_6 : _GEN_821; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_823 = 5'h7 == upperNodeIndex[4:0] ? frequency_7 : _GEN_822; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_824 = 5'h8 == upperNodeIndex[4:0] ? frequency_8 : _GEN_823; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_825 = 5'h9 == upperNodeIndex[4:0] ? frequency_9 : _GEN_824; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_826 = 5'ha == upperNodeIndex[4:0] ? frequency_10 : _GEN_825; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_827 = 5'hb == upperNodeIndex[4:0] ? frequency_11 : _GEN_826; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_828 = 5'hc == upperNodeIndex[4:0] ? frequency_12 : _GEN_827; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_829 = 5'hd == upperNodeIndex[4:0] ? frequency_13 : _GEN_828; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_830 = 5'he == upperNodeIndex[4:0] ? frequency_14 : _GEN_829; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_831 = 5'hf == upperNodeIndex[4:0] ? frequency_15 : _GEN_830; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_832 = 5'h10 == upperNodeIndex[4:0] ? frequency_16 : _GEN_831; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_833 = 5'h11 == upperNodeIndex[4:0] ? frequency_17 : _GEN_832; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_834 = 5'h12 == upperNodeIndex[4:0] ? frequency_18 : _GEN_833; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_835 = 5'h13 == upperNodeIndex[4:0] ? frequency_19 : _GEN_834; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_836 = 5'h14 == upperNodeIndex[4:0] ? frequency_20 : _GEN_835; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_837 = 5'h15 == upperNodeIndex[4:0] ? frequency_21 : _GEN_836; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_838 = 5'h16 == upperNodeIndex[4:0] ? frequency_22 : _GEN_837; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_839 = 5'h17 == upperNodeIndex[4:0] ? frequency_23 : _GEN_838; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_840 = 5'h18 == upperNodeIndex[4:0] ? frequency_24 : _GEN_839; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_841 = 5'h19 == upperNodeIndex[4:0] ? frequency_25 : _GEN_840; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_842 = 5'h1a == upperNodeIndex[4:0] ? frequency_26 : _GEN_841; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_843 = 5'h1b == upperNodeIndex[4:0] ? frequency_27 : _GEN_842; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_844 = 5'h1c == upperNodeIndex[4:0] ? frequency_28 : _GEN_843; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_845 = 5'h1d == upperNodeIndex[4:0] ? frequency_29 : _GEN_844; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_846 = 5'h1e == upperNodeIndex[4:0] ? frequency_30 : _GEN_845; // @[treeGenerator.scala 152:62]
  wire [12:0] _GEN_847 = 5'h1f == upperNodeIndex[4:0] ? frequency_31 : _GEN_846; // @[treeGenerator.scala 152:62]
  wire  _T_320 = newFrequency == _GEN_847; // @[treeGenerator.scala 152:62]
  wire  _T_321 = _T_318 | _T_320; // @[treeGenerator.scala 152:45]
  wire [12:0] _GEN_849 = 5'h1 == lowerNodeIndex[4:0] ? frequency_1 : frequency_0; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_850 = 5'h2 == lowerNodeIndex[4:0] ? frequency_2 : _GEN_849; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_851 = 5'h3 == lowerNodeIndex[4:0] ? frequency_3 : _GEN_850; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_852 = 5'h4 == lowerNodeIndex[4:0] ? frequency_4 : _GEN_851; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_853 = 5'h5 == lowerNodeIndex[4:0] ? frequency_5 : _GEN_852; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_854 = 5'h6 == lowerNodeIndex[4:0] ? frequency_6 : _GEN_853; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_855 = 5'h7 == lowerNodeIndex[4:0] ? frequency_7 : _GEN_854; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_856 = 5'h8 == lowerNodeIndex[4:0] ? frequency_8 : _GEN_855; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_857 = 5'h9 == lowerNodeIndex[4:0] ? frequency_9 : _GEN_856; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_858 = 5'ha == lowerNodeIndex[4:0] ? frequency_10 : _GEN_857; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_859 = 5'hb == lowerNodeIndex[4:0] ? frequency_11 : _GEN_858; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_860 = 5'hc == lowerNodeIndex[4:0] ? frequency_12 : _GEN_859; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_861 = 5'hd == lowerNodeIndex[4:0] ? frequency_13 : _GEN_860; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_862 = 5'he == lowerNodeIndex[4:0] ? frequency_14 : _GEN_861; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_863 = 5'hf == lowerNodeIndex[4:0] ? frequency_15 : _GEN_862; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_864 = 5'h10 == lowerNodeIndex[4:0] ? frequency_16 : _GEN_863; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_865 = 5'h11 == lowerNodeIndex[4:0] ? frequency_17 : _GEN_864; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_866 = 5'h12 == lowerNodeIndex[4:0] ? frequency_18 : _GEN_865; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_867 = 5'h13 == lowerNodeIndex[4:0] ? frequency_19 : _GEN_866; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_868 = 5'h14 == lowerNodeIndex[4:0] ? frequency_20 : _GEN_867; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_869 = 5'h15 == lowerNodeIndex[4:0] ? frequency_21 : _GEN_868; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_870 = 5'h16 == lowerNodeIndex[4:0] ? frequency_22 : _GEN_869; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_871 = 5'h17 == lowerNodeIndex[4:0] ? frequency_23 : _GEN_870; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_872 = 5'h18 == lowerNodeIndex[4:0] ? frequency_24 : _GEN_871; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_873 = 5'h19 == lowerNodeIndex[4:0] ? frequency_25 : _GEN_872; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_874 = 5'h1a == lowerNodeIndex[4:0] ? frequency_26 : _GEN_873; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_875 = 5'h1b == lowerNodeIndex[4:0] ? frequency_27 : _GEN_874; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_876 = 5'h1c == lowerNodeIndex[4:0] ? frequency_28 : _GEN_875; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_877 = 5'h1d == lowerNodeIndex[4:0] ? frequency_29 : _GEN_876; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_878 = 5'h1e == lowerNodeIndex[4:0] ? frequency_30 : _GEN_877; // @[treeGenerator.scala 159:36]
  wire [12:0] _GEN_879 = 5'h1f == lowerNodeIndex[4:0] ? frequency_31 : _GEN_878; // @[treeGenerator.scala 159:36]
  wire  _T_323 = _GEN_879 == newFrequency; // @[treeGenerator.scala 159:36]
  wire  _T_325 = _GEN_847 > newFrequency; // @[treeGenerator.scala 160:40]
  wire  _T_327 = _GEN_879 < newFrequency; // @[treeGenerator.scala 162:13]
  wire  _T_328 = _T_325 & _T_327; // @[treeGenerator.scala 160:56]
  wire [5:0] _T_330 = upperNodeIndex + 6'h1; // @[treeGenerator.scala 162:50]
  wire  _T_331 = _T_330 == lowerNodeIndex; // @[treeGenerator.scala 162:57]
  wire  _T_332 = _T_328 & _T_331; // @[treeGenerator.scala 162:30]
  wire  _T_333 = _T_323 | _T_332; // @[treeGenerator.scala 159:54]
  wire [5:0] _GEN_945 = _T_333 ? lowerNodeIndex : 6'h0; // @[treeGenerator.scala 163:9]
  wire  _GEN_946 = _T_321 | _T_333; // @[treeGenerator.scala 155:9]
  wire [5:0] _GEN_947 = _T_321 ? upperNodeIndex : _GEN_945; // @[treeGenerator.scala 155:9]
  wire [5:0] _GEN_1271 = _T_317 ? _GEN_947 : 6'h0; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_1636 = _T_284 ? 6'h0 : _GEN_1271; // @[Conditional.scala 39:67]
  wire [5:0] matchedIndex = _T_32 ? 6'h0 : _GEN_1636; // @[Conditional.scala 40:58]
  wire  _T_334 = 6'h0 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_336 = 6'h1 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_337 = 6'h1 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_338 = 6'h2 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_339 = 6'h2 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_340 = 6'h3 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_341 = 6'h3 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_342 = 6'h4 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_343 = 6'h4 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_344 = 6'h5 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_345 = 6'h5 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_346 = 6'h6 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_347 = 6'h6 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_348 = 6'h7 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_349 = 6'h7 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_350 = 6'h8 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_351 = 6'h8 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_352 = 6'h9 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_353 = 6'h9 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_354 = 6'ha == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_355 = 6'ha > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_356 = 6'hb == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_357 = 6'hb > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_358 = 6'hc == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_359 = 6'hc > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_360 = 6'hd == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_361 = 6'hd > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_362 = 6'he == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_363 = 6'he > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_364 = 6'hf == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_365 = 6'hf > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_366 = 6'h10 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_367 = 6'h10 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_368 = 6'h11 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_369 = 6'h11 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_370 = 6'h12 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_371 = 6'h12 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_372 = 6'h13 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_373 = 6'h13 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_374 = 6'h14 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_375 = 6'h14 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_376 = 6'h15 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_377 = 6'h15 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_378 = 6'h16 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_379 = 6'h16 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_380 = 6'h17 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_381 = 6'h17 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_382 = 6'h18 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_383 = 6'h18 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_384 = 6'h19 == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_385 = 6'h19 > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_386 = 6'h1a == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_387 = 6'h1a > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_388 = 6'h1b == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_389 = 6'h1b > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_390 = 6'h1c == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_391 = 6'h1c > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_392 = 6'h1d == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_393 = 6'h1d > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_394 = 6'h1e == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_395 = 6'h1e > matchedIndex; // @[treeGenerator.scala 176:30]
  wire  _T_396 = 6'h1f == matchedIndex; // @[treeGenerator.scala 172:24]
  wire  _T_397 = 6'h1f > matchedIndex; // @[treeGenerator.scala 176:30]
  wire [5:0] _T_399 = lowerNodeIndex - upperNodeIndex; // @[treeGenerator.scala 185:37]
  wire [5:0] _T_400 = _T_399 / 6'h2; // @[treeGenerator.scala 185:55]
  wire [5:0] _T_402 = _T_400 + upperNodeIndex; // @[treeGenerator.scala 185:61]
  wire [12:0] _GEN_1138 = 5'h1 == _T_402[4:0] ? frequency_1 : frequency_0; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1139 = 5'h2 == _T_402[4:0] ? frequency_2 : _GEN_1138; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1140 = 5'h3 == _T_402[4:0] ? frequency_3 : _GEN_1139; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1141 = 5'h4 == _T_402[4:0] ? frequency_4 : _GEN_1140; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1142 = 5'h5 == _T_402[4:0] ? frequency_5 : _GEN_1141; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1143 = 5'h6 == _T_402[4:0] ? frequency_6 : _GEN_1142; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1144 = 5'h7 == _T_402[4:0] ? frequency_7 : _GEN_1143; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1145 = 5'h8 == _T_402[4:0] ? frequency_8 : _GEN_1144; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1146 = 5'h9 == _T_402[4:0] ? frequency_9 : _GEN_1145; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1147 = 5'ha == _T_402[4:0] ? frequency_10 : _GEN_1146; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1148 = 5'hb == _T_402[4:0] ? frequency_11 : _GEN_1147; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1149 = 5'hc == _T_402[4:0] ? frequency_12 : _GEN_1148; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1150 = 5'hd == _T_402[4:0] ? frequency_13 : _GEN_1149; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1151 = 5'he == _T_402[4:0] ? frequency_14 : _GEN_1150; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1152 = 5'hf == _T_402[4:0] ? frequency_15 : _GEN_1151; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1153 = 5'h10 == _T_402[4:0] ? frequency_16 : _GEN_1152; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1154 = 5'h11 == _T_402[4:0] ? frequency_17 : _GEN_1153; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1155 = 5'h12 == _T_402[4:0] ? frequency_18 : _GEN_1154; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1156 = 5'h13 == _T_402[4:0] ? frequency_19 : _GEN_1155; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1157 = 5'h14 == _T_402[4:0] ? frequency_20 : _GEN_1156; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1158 = 5'h15 == _T_402[4:0] ? frequency_21 : _GEN_1157; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1159 = 5'h16 == _T_402[4:0] ? frequency_22 : _GEN_1158; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1160 = 5'h17 == _T_402[4:0] ? frequency_23 : _GEN_1159; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1161 = 5'h18 == _T_402[4:0] ? frequency_24 : _GEN_1160; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1162 = 5'h19 == _T_402[4:0] ? frequency_25 : _GEN_1161; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1163 = 5'h1a == _T_402[4:0] ? frequency_26 : _GEN_1162; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1164 = 5'h1b == _T_402[4:0] ? frequency_27 : _GEN_1163; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1165 = 5'h1c == _T_402[4:0] ? frequency_28 : _GEN_1164; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1166 = 5'h1d == _T_402[4:0] ? frequency_29 : _GEN_1165; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1167 = 5'h1e == _T_402[4:0] ? frequency_30 : _GEN_1166; // @[treeGenerator.scala 185:79]
  wire [12:0] _GEN_1168 = 5'h1f == _T_402[4:0] ? frequency_31 : _GEN_1167; // @[treeGenerator.scala 185:79]
  wire  _T_404 = _GEN_1168 < newFrequency; // @[treeGenerator.scala 185:79]
  wire  _GEN_1270 = _T_317 & _GEN_946; // @[Conditional.scala 39:67]
  wire  _GEN_1635 = _T_284 ? 1'h0 : _GEN_1270; // @[Conditional.scala 39:67]
  wire  searchCompleted = _T_32 ? 1'h0 : _GEN_1635; // @[Conditional.scala 40:58]
  assign io_outputs_leftNode_0 = leftNode_0; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_1 = leftNode_1; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_2 = leftNode_2; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_3 = leftNode_3; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_4 = leftNode_4; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_5 = leftNode_5; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_6 = leftNode_6; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_7 = leftNode_7; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_8 = leftNode_8; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_9 = leftNode_9; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_10 = leftNode_10; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_11 = leftNode_11; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_12 = leftNode_12; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_13 = leftNode_13; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_14 = leftNode_14; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_15 = leftNode_15; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_16 = leftNode_16; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_17 = leftNode_17; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_18 = leftNode_18; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_19 = leftNode_19; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_20 = leftNode_20; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_21 = leftNode_21; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_22 = leftNode_22; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_23 = leftNode_23; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_24 = leftNode_24; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_25 = leftNode_25; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_26 = leftNode_26; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_27 = leftNode_27; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_28 = leftNode_28; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_29 = leftNode_29; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_30 = leftNode_30; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_31 = leftNode_31; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_32 = leftNode_32; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_33 = leftNode_33; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_34 = leftNode_34; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_35 = leftNode_35; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_36 = leftNode_36; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_37 = leftNode_37; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_38 = leftNode_38; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_39 = leftNode_39; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_40 = leftNode_40; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_41 = leftNode_41; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_42 = leftNode_42; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_43 = leftNode_43; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_44 = leftNode_44; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_45 = leftNode_45; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_46 = leftNode_46; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_47 = leftNode_47; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_48 = leftNode_48; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_49 = leftNode_49; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_50 = leftNode_50; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_51 = leftNode_51; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_52 = leftNode_52; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_53 = leftNode_53; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_54 = leftNode_54; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_55 = leftNode_55; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_56 = leftNode_56; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_57 = leftNode_57; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_58 = leftNode_58; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_59 = leftNode_59; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_60 = leftNode_60; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_61 = leftNode_61; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_62 = leftNode_62; // @[treeGenerator.scala 195:23]
  assign io_outputs_leftNode_63 = leftNode_63; // @[treeGenerator.scala 195:23]
  assign io_outputs_rightNode_0 = rightNode_0; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_1 = rightNode_1; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_2 = rightNode_2; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_3 = rightNode_3; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_4 = rightNode_4; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_5 = rightNode_5; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_6 = rightNode_6; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_7 = rightNode_7; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_8 = rightNode_8; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_9 = rightNode_9; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_10 = rightNode_10; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_11 = rightNode_11; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_12 = rightNode_12; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_13 = rightNode_13; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_14 = rightNode_14; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_15 = rightNode_15; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_16 = rightNode_16; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_17 = rightNode_17; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_18 = rightNode_18; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_19 = rightNode_19; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_20 = rightNode_20; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_21 = rightNode_21; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_22 = rightNode_22; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_23 = rightNode_23; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_24 = rightNode_24; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_25 = rightNode_25; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_26 = rightNode_26; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_27 = rightNode_27; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_28 = rightNode_28; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_29 = rightNode_29; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_30 = rightNode_30; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_31 = rightNode_31; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_32 = rightNode_32; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_33 = rightNode_33; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_34 = rightNode_34; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_35 = rightNode_35; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_36 = rightNode_36; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_37 = rightNode_37; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_38 = rightNode_38; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_39 = rightNode_39; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_40 = rightNode_40; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_41 = rightNode_41; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_42 = rightNode_42; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_43 = rightNode_43; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_44 = rightNode_44; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_45 = rightNode_45; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_46 = rightNode_46; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_47 = rightNode_47; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_48 = rightNode_48; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_49 = rightNode_49; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_50 = rightNode_50; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_51 = rightNode_51; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_52 = rightNode_52; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_53 = rightNode_53; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_54 = rightNode_54; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_55 = rightNode_55; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_56 = rightNode_56; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_57 = rightNode_57; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_58 = rightNode_58; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_59 = rightNode_59; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_60 = rightNode_60; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_61 = rightNode_61; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_62 = rightNode_62; // @[treeGenerator.scala 196:24]
  assign io_outputs_rightNode_63 = rightNode_63; // @[treeGenerator.scala 196:24]
  assign io_outputs_leftNodeIsCharacter_0 = leftNodeIsCharacter_0; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_1 = leftNodeIsCharacter_1; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_2 = leftNodeIsCharacter_2; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_3 = leftNodeIsCharacter_3; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_4 = leftNodeIsCharacter_4; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_5 = leftNodeIsCharacter_5; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_6 = leftNodeIsCharacter_6; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_7 = leftNodeIsCharacter_7; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_8 = leftNodeIsCharacter_8; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_9 = leftNodeIsCharacter_9; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_10 = leftNodeIsCharacter_10; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_11 = leftNodeIsCharacter_11; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_12 = leftNodeIsCharacter_12; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_13 = leftNodeIsCharacter_13; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_14 = leftNodeIsCharacter_14; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_15 = leftNodeIsCharacter_15; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_16 = leftNodeIsCharacter_16; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_17 = leftNodeIsCharacter_17; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_18 = leftNodeIsCharacter_18; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_19 = leftNodeIsCharacter_19; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_20 = leftNodeIsCharacter_20; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_21 = leftNodeIsCharacter_21; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_22 = leftNodeIsCharacter_22; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_23 = leftNodeIsCharacter_23; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_24 = leftNodeIsCharacter_24; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_25 = leftNodeIsCharacter_25; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_26 = leftNodeIsCharacter_26; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_27 = leftNodeIsCharacter_27; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_28 = leftNodeIsCharacter_28; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_29 = leftNodeIsCharacter_29; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_30 = leftNodeIsCharacter_30; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_31 = leftNodeIsCharacter_31; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_32 = leftNodeIsCharacter_32; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_33 = leftNodeIsCharacter_33; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_34 = leftNodeIsCharacter_34; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_35 = leftNodeIsCharacter_35; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_36 = leftNodeIsCharacter_36; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_37 = leftNodeIsCharacter_37; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_38 = leftNodeIsCharacter_38; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_39 = leftNodeIsCharacter_39; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_40 = leftNodeIsCharacter_40; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_41 = leftNodeIsCharacter_41; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_42 = leftNodeIsCharacter_42; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_43 = leftNodeIsCharacter_43; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_44 = leftNodeIsCharacter_44; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_45 = leftNodeIsCharacter_45; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_46 = leftNodeIsCharacter_46; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_47 = leftNodeIsCharacter_47; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_48 = leftNodeIsCharacter_48; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_49 = leftNodeIsCharacter_49; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_50 = leftNodeIsCharacter_50; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_51 = leftNodeIsCharacter_51; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_52 = leftNodeIsCharacter_52; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_53 = leftNodeIsCharacter_53; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_54 = leftNodeIsCharacter_54; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_55 = leftNodeIsCharacter_55; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_56 = leftNodeIsCharacter_56; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_57 = leftNodeIsCharacter_57; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_58 = leftNodeIsCharacter_58; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_59 = leftNodeIsCharacter_59; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_60 = leftNodeIsCharacter_60; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_61 = leftNodeIsCharacter_61; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_62 = leftNodeIsCharacter_62; // @[treeGenerator.scala 197:34]
  assign io_outputs_leftNodeIsCharacter_63 = leftNodeIsCharacter_63; // @[treeGenerator.scala 197:34]
  assign io_outputs_rightNodeIsCharacter_0 = rightNodeIsCharacter_0; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_1 = rightNodeIsCharacter_1; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_2 = rightNodeIsCharacter_2; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_3 = rightNodeIsCharacter_3; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_4 = rightNodeIsCharacter_4; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_5 = rightNodeIsCharacter_5; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_6 = rightNodeIsCharacter_6; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_7 = rightNodeIsCharacter_7; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_8 = rightNodeIsCharacter_8; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_9 = rightNodeIsCharacter_9; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_10 = rightNodeIsCharacter_10; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_11 = rightNodeIsCharacter_11; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_12 = rightNodeIsCharacter_12; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_13 = rightNodeIsCharacter_13; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_14 = rightNodeIsCharacter_14; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_15 = rightNodeIsCharacter_15; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_16 = rightNodeIsCharacter_16; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_17 = rightNodeIsCharacter_17; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_18 = rightNodeIsCharacter_18; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_19 = rightNodeIsCharacter_19; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_20 = rightNodeIsCharacter_20; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_21 = rightNodeIsCharacter_21; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_22 = rightNodeIsCharacter_22; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_23 = rightNodeIsCharacter_23; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_24 = rightNodeIsCharacter_24; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_25 = rightNodeIsCharacter_25; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_26 = rightNodeIsCharacter_26; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_27 = rightNodeIsCharacter_27; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_28 = rightNodeIsCharacter_28; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_29 = rightNodeIsCharacter_29; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_30 = rightNodeIsCharacter_30; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_31 = rightNodeIsCharacter_31; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_32 = rightNodeIsCharacter_32; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_33 = rightNodeIsCharacter_33; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_34 = rightNodeIsCharacter_34; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_35 = rightNodeIsCharacter_35; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_36 = rightNodeIsCharacter_36; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_37 = rightNodeIsCharacter_37; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_38 = rightNodeIsCharacter_38; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_39 = rightNodeIsCharacter_39; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_40 = rightNodeIsCharacter_40; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_41 = rightNodeIsCharacter_41; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_42 = rightNodeIsCharacter_42; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_43 = rightNodeIsCharacter_43; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_44 = rightNodeIsCharacter_44; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_45 = rightNodeIsCharacter_45; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_46 = rightNodeIsCharacter_46; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_47 = rightNodeIsCharacter_47; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_48 = rightNodeIsCharacter_48; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_49 = rightNodeIsCharacter_49; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_50 = rightNodeIsCharacter_50; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_51 = rightNodeIsCharacter_51; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_52 = rightNodeIsCharacter_52; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_53 = rightNodeIsCharacter_53; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_54 = rightNodeIsCharacter_54; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_55 = rightNodeIsCharacter_55; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_56 = rightNodeIsCharacter_56; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_57 = rightNodeIsCharacter_57; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_58 = rightNodeIsCharacter_58; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_59 = rightNodeIsCharacter_59; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_60 = rightNodeIsCharacter_60; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_61 = rightNodeIsCharacter_61; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_62 = rightNodeIsCharacter_62; // @[treeGenerator.scala 198:35]
  assign io_outputs_rightNodeIsCharacter_63 = rightNodeIsCharacter_63; // @[treeGenerator.scala 198:35]
  assign io_outputs_validNodes = validNodes; // @[treeGenerator.scala 199:25]
  assign io_outputs_validCharacters = validCharacters; // @[treeGenerator.scala 200:30]
  assign io_finished = state == 2'h0; // @[treeGenerator.scala 201:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  frequency_0 = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  frequency_1 = _RAND_1[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  frequency_2 = _RAND_2[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  frequency_3 = _RAND_3[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  frequency_4 = _RAND_4[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  frequency_5 = _RAND_5[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  frequency_6 = _RAND_6[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  frequency_7 = _RAND_7[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  frequency_8 = _RAND_8[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  frequency_9 = _RAND_9[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  frequency_10 = _RAND_10[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  frequency_11 = _RAND_11[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  frequency_12 = _RAND_12[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  frequency_13 = _RAND_13[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  frequency_14 = _RAND_14[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  frequency_15 = _RAND_15[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  frequency_16 = _RAND_16[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  frequency_17 = _RAND_17[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  frequency_18 = _RAND_18[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  frequency_19 = _RAND_19[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  frequency_20 = _RAND_20[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  frequency_21 = _RAND_21[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  frequency_22 = _RAND_22[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  frequency_23 = _RAND_23[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  frequency_24 = _RAND_24[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  frequency_25 = _RAND_25[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  frequency_26 = _RAND_26[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  frequency_27 = _RAND_27[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  frequency_28 = _RAND_28[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  frequency_29 = _RAND_29[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  frequency_30 = _RAND_30[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  frequency_31 = _RAND_31[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  pointerOrCharacter_0 = _RAND_32[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  pointerOrCharacter_1 = _RAND_33[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  pointerOrCharacter_2 = _RAND_34[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  pointerOrCharacter_3 = _RAND_35[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  pointerOrCharacter_4 = _RAND_36[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  pointerOrCharacter_5 = _RAND_37[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  pointerOrCharacter_6 = _RAND_38[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  pointerOrCharacter_7 = _RAND_39[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  pointerOrCharacter_8 = _RAND_40[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  pointerOrCharacter_9 = _RAND_41[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  pointerOrCharacter_10 = _RAND_42[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  pointerOrCharacter_11 = _RAND_43[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  pointerOrCharacter_12 = _RAND_44[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  pointerOrCharacter_13 = _RAND_45[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  pointerOrCharacter_14 = _RAND_46[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  pointerOrCharacter_15 = _RAND_47[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  pointerOrCharacter_16 = _RAND_48[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  pointerOrCharacter_17 = _RAND_49[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  pointerOrCharacter_18 = _RAND_50[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  pointerOrCharacter_19 = _RAND_51[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  pointerOrCharacter_20 = _RAND_52[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  pointerOrCharacter_21 = _RAND_53[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  pointerOrCharacter_22 = _RAND_54[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  pointerOrCharacter_23 = _RAND_55[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  pointerOrCharacter_24 = _RAND_56[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  pointerOrCharacter_25 = _RAND_57[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  pointerOrCharacter_26 = _RAND_58[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  pointerOrCharacter_27 = _RAND_59[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  pointerOrCharacter_28 = _RAND_60[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  pointerOrCharacter_29 = _RAND_61[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  pointerOrCharacter_30 = _RAND_62[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  pointerOrCharacter_31 = _RAND_63[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  isCharacter_0 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  isCharacter_1 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  isCharacter_2 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  isCharacter_3 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  isCharacter_4 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  isCharacter_5 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  isCharacter_6 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  isCharacter_7 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  isCharacter_8 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  isCharacter_9 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  isCharacter_10 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  isCharacter_11 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  isCharacter_12 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  isCharacter_13 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  isCharacter_14 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  isCharacter_15 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  isCharacter_16 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  isCharacter_17 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  isCharacter_18 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  isCharacter_19 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  isCharacter_20 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  isCharacter_21 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  isCharacter_22 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  isCharacter_23 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  isCharacter_24 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  isCharacter_25 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  isCharacter_26 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  isCharacter_27 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  isCharacter_28 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  isCharacter_29 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  isCharacter_30 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  isCharacter_31 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  newFrequency = _RAND_96[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  newPointer = _RAND_97[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  validRoots = _RAND_98[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  leftNode_0 = _RAND_99[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  leftNode_1 = _RAND_100[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  leftNode_2 = _RAND_101[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  leftNode_3 = _RAND_102[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  leftNode_4 = _RAND_103[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  leftNode_5 = _RAND_104[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  leftNode_6 = _RAND_105[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  leftNode_7 = _RAND_106[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  leftNode_8 = _RAND_107[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  leftNode_9 = _RAND_108[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  leftNode_10 = _RAND_109[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  leftNode_11 = _RAND_110[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  leftNode_12 = _RAND_111[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  leftNode_13 = _RAND_112[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  leftNode_14 = _RAND_113[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  leftNode_15 = _RAND_114[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  leftNode_16 = _RAND_115[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  leftNode_17 = _RAND_116[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  leftNode_18 = _RAND_117[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  leftNode_19 = _RAND_118[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  leftNode_20 = _RAND_119[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  leftNode_21 = _RAND_120[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  leftNode_22 = _RAND_121[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  leftNode_23 = _RAND_122[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  leftNode_24 = _RAND_123[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  leftNode_25 = _RAND_124[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  leftNode_26 = _RAND_125[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  leftNode_27 = _RAND_126[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  leftNode_28 = _RAND_127[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  leftNode_29 = _RAND_128[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  leftNode_30 = _RAND_129[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  leftNode_31 = _RAND_130[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  leftNode_32 = _RAND_131[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  leftNode_33 = _RAND_132[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  leftNode_34 = _RAND_133[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  leftNode_35 = _RAND_134[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  leftNode_36 = _RAND_135[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  leftNode_37 = _RAND_136[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  leftNode_38 = _RAND_137[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  leftNode_39 = _RAND_138[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  leftNode_40 = _RAND_139[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  leftNode_41 = _RAND_140[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  leftNode_42 = _RAND_141[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  leftNode_43 = _RAND_142[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  leftNode_44 = _RAND_143[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  leftNode_45 = _RAND_144[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  leftNode_46 = _RAND_145[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  leftNode_47 = _RAND_146[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  leftNode_48 = _RAND_147[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  leftNode_49 = _RAND_148[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  leftNode_50 = _RAND_149[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  leftNode_51 = _RAND_150[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  leftNode_52 = _RAND_151[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  leftNode_53 = _RAND_152[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  leftNode_54 = _RAND_153[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  leftNode_55 = _RAND_154[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  leftNode_56 = _RAND_155[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  leftNode_57 = _RAND_156[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  leftNode_58 = _RAND_157[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  leftNode_59 = _RAND_158[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  leftNode_60 = _RAND_159[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  leftNode_61 = _RAND_160[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  leftNode_62 = _RAND_161[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  leftNode_63 = _RAND_162[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  rightNode_0 = _RAND_163[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  rightNode_1 = _RAND_164[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  rightNode_2 = _RAND_165[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  rightNode_3 = _RAND_166[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  rightNode_4 = _RAND_167[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  rightNode_5 = _RAND_168[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  rightNode_6 = _RAND_169[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  rightNode_7 = _RAND_170[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  rightNode_8 = _RAND_171[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  rightNode_9 = _RAND_172[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  rightNode_10 = _RAND_173[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  rightNode_11 = _RAND_174[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  rightNode_12 = _RAND_175[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  rightNode_13 = _RAND_176[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  rightNode_14 = _RAND_177[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  rightNode_15 = _RAND_178[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  rightNode_16 = _RAND_179[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  rightNode_17 = _RAND_180[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  rightNode_18 = _RAND_181[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  rightNode_19 = _RAND_182[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  rightNode_20 = _RAND_183[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  rightNode_21 = _RAND_184[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  rightNode_22 = _RAND_185[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  rightNode_23 = _RAND_186[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  rightNode_24 = _RAND_187[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  rightNode_25 = _RAND_188[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  rightNode_26 = _RAND_189[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  rightNode_27 = _RAND_190[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  rightNode_28 = _RAND_191[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  rightNode_29 = _RAND_192[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  rightNode_30 = _RAND_193[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  rightNode_31 = _RAND_194[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  rightNode_32 = _RAND_195[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  rightNode_33 = _RAND_196[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  rightNode_34 = _RAND_197[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  rightNode_35 = _RAND_198[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  rightNode_36 = _RAND_199[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  rightNode_37 = _RAND_200[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  rightNode_38 = _RAND_201[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  rightNode_39 = _RAND_202[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  rightNode_40 = _RAND_203[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  rightNode_41 = _RAND_204[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  rightNode_42 = _RAND_205[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  rightNode_43 = _RAND_206[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  rightNode_44 = _RAND_207[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  rightNode_45 = _RAND_208[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  rightNode_46 = _RAND_209[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  rightNode_47 = _RAND_210[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  rightNode_48 = _RAND_211[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  rightNode_49 = _RAND_212[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  rightNode_50 = _RAND_213[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  rightNode_51 = _RAND_214[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  rightNode_52 = _RAND_215[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  rightNode_53 = _RAND_216[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  rightNode_54 = _RAND_217[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  rightNode_55 = _RAND_218[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  rightNode_56 = _RAND_219[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  rightNode_57 = _RAND_220[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  rightNode_58 = _RAND_221[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  rightNode_59 = _RAND_222[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  rightNode_60 = _RAND_223[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  rightNode_61 = _RAND_224[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  rightNode_62 = _RAND_225[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  rightNode_63 = _RAND_226[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  leftNodeIsCharacter_0 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  leftNodeIsCharacter_1 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  leftNodeIsCharacter_2 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  leftNodeIsCharacter_3 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  leftNodeIsCharacter_4 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  leftNodeIsCharacter_5 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  leftNodeIsCharacter_6 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  leftNodeIsCharacter_7 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  leftNodeIsCharacter_8 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  leftNodeIsCharacter_9 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  leftNodeIsCharacter_10 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  leftNodeIsCharacter_11 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  leftNodeIsCharacter_12 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  leftNodeIsCharacter_13 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  leftNodeIsCharacter_14 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  leftNodeIsCharacter_15 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  leftNodeIsCharacter_16 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  leftNodeIsCharacter_17 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  leftNodeIsCharacter_18 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  leftNodeIsCharacter_19 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  leftNodeIsCharacter_20 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  leftNodeIsCharacter_21 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  leftNodeIsCharacter_22 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  leftNodeIsCharacter_23 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  leftNodeIsCharacter_24 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  leftNodeIsCharacter_25 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  leftNodeIsCharacter_26 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  leftNodeIsCharacter_27 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  leftNodeIsCharacter_28 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  leftNodeIsCharacter_29 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  leftNodeIsCharacter_30 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  leftNodeIsCharacter_31 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  leftNodeIsCharacter_32 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  leftNodeIsCharacter_33 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  leftNodeIsCharacter_34 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  leftNodeIsCharacter_35 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  leftNodeIsCharacter_36 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  leftNodeIsCharacter_37 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  leftNodeIsCharacter_38 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  leftNodeIsCharacter_39 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  leftNodeIsCharacter_40 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  leftNodeIsCharacter_41 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  leftNodeIsCharacter_42 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  leftNodeIsCharacter_43 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  leftNodeIsCharacter_44 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  leftNodeIsCharacter_45 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  leftNodeIsCharacter_46 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  leftNodeIsCharacter_47 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  leftNodeIsCharacter_48 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  leftNodeIsCharacter_49 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  leftNodeIsCharacter_50 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  leftNodeIsCharacter_51 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  leftNodeIsCharacter_52 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  leftNodeIsCharacter_53 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  leftNodeIsCharacter_54 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  leftNodeIsCharacter_55 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  leftNodeIsCharacter_56 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  leftNodeIsCharacter_57 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  leftNodeIsCharacter_58 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  leftNodeIsCharacter_59 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  leftNodeIsCharacter_60 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  leftNodeIsCharacter_61 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  leftNodeIsCharacter_62 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  leftNodeIsCharacter_63 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  rightNodeIsCharacter_0 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  rightNodeIsCharacter_1 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  rightNodeIsCharacter_2 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  rightNodeIsCharacter_3 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  rightNodeIsCharacter_4 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  rightNodeIsCharacter_5 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  rightNodeIsCharacter_6 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  rightNodeIsCharacter_7 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  rightNodeIsCharacter_8 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  rightNodeIsCharacter_9 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  rightNodeIsCharacter_10 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  rightNodeIsCharacter_11 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  rightNodeIsCharacter_12 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  rightNodeIsCharacter_13 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  rightNodeIsCharacter_14 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  rightNodeIsCharacter_15 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  rightNodeIsCharacter_16 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  rightNodeIsCharacter_17 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  rightNodeIsCharacter_18 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  rightNodeIsCharacter_19 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  rightNodeIsCharacter_20 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  rightNodeIsCharacter_21 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  rightNodeIsCharacter_22 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  rightNodeIsCharacter_23 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  rightNodeIsCharacter_24 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  rightNodeIsCharacter_25 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  rightNodeIsCharacter_26 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  rightNodeIsCharacter_27 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  rightNodeIsCharacter_28 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  rightNodeIsCharacter_29 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  rightNodeIsCharacter_30 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  rightNodeIsCharacter_31 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  rightNodeIsCharacter_32 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  rightNodeIsCharacter_33 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  rightNodeIsCharacter_34 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  rightNodeIsCharacter_35 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  rightNodeIsCharacter_36 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  rightNodeIsCharacter_37 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  rightNodeIsCharacter_38 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  rightNodeIsCharacter_39 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  rightNodeIsCharacter_40 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  rightNodeIsCharacter_41 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  rightNodeIsCharacter_42 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  rightNodeIsCharacter_43 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  rightNodeIsCharacter_44 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  rightNodeIsCharacter_45 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  rightNodeIsCharacter_46 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  rightNodeIsCharacter_47 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  rightNodeIsCharacter_48 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  rightNodeIsCharacter_49 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  rightNodeIsCharacter_50 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  rightNodeIsCharacter_51 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  rightNodeIsCharacter_52 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  rightNodeIsCharacter_53 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  rightNodeIsCharacter_54 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  rightNodeIsCharacter_55 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  rightNodeIsCharacter_56 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  rightNodeIsCharacter_57 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  rightNodeIsCharacter_58 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  rightNodeIsCharacter_59 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  rightNodeIsCharacter_60 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  rightNodeIsCharacter_61 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  rightNodeIsCharacter_62 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  rightNodeIsCharacter_63 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  upperNodeIndex = _RAND_355[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  lowerNodeIndex = _RAND_356[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  validNodes = _RAND_357[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  validCharacters = _RAND_358[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  state = _RAND_359[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_32) begin
      if (io_start) begin
        frequency_0 <= io_inputs_sortedFrequency_0;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_334) begin
            frequency_0 <= newFrequency;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_1 <= io_inputs_sortedFrequency_1;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_336) begin
            frequency_1 <= newFrequency;
          end else if (_T_337) begin
            frequency_1 <= frequency_0;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_2 <= io_inputs_sortedFrequency_2;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_338) begin
            frequency_2 <= newFrequency;
          end else if (_T_339) begin
            frequency_2 <= frequency_1;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_3 <= io_inputs_sortedFrequency_3;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_340) begin
            frequency_3 <= newFrequency;
          end else if (_T_341) begin
            frequency_3 <= frequency_2;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_4 <= io_inputs_sortedFrequency_4;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_342) begin
            frequency_4 <= newFrequency;
          end else if (_T_343) begin
            frequency_4 <= frequency_3;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_5 <= io_inputs_sortedFrequency_5;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_344) begin
            frequency_5 <= newFrequency;
          end else if (_T_345) begin
            frequency_5 <= frequency_4;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_6 <= io_inputs_sortedFrequency_6;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_346) begin
            frequency_6 <= newFrequency;
          end else if (_T_347) begin
            frequency_6 <= frequency_5;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_7 <= io_inputs_sortedFrequency_7;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_348) begin
            frequency_7 <= newFrequency;
          end else if (_T_349) begin
            frequency_7 <= frequency_6;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_8 <= io_inputs_sortedFrequency_8;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_350) begin
            frequency_8 <= newFrequency;
          end else if (_T_351) begin
            frequency_8 <= frequency_7;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_9 <= io_inputs_sortedFrequency_9;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_352) begin
            frequency_9 <= newFrequency;
          end else if (_T_353) begin
            frequency_9 <= frequency_8;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_10 <= io_inputs_sortedFrequency_10;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_354) begin
            frequency_10 <= newFrequency;
          end else if (_T_355) begin
            frequency_10 <= frequency_9;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_11 <= io_inputs_sortedFrequency_11;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_356) begin
            frequency_11 <= newFrequency;
          end else if (_T_357) begin
            frequency_11 <= frequency_10;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_12 <= io_inputs_sortedFrequency_12;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_358) begin
            frequency_12 <= newFrequency;
          end else if (_T_359) begin
            frequency_12 <= frequency_11;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_13 <= io_inputs_sortedFrequency_13;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_360) begin
            frequency_13 <= newFrequency;
          end else if (_T_361) begin
            frequency_13 <= frequency_12;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_14 <= io_inputs_sortedFrequency_14;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_362) begin
            frequency_14 <= newFrequency;
          end else if (_T_363) begin
            frequency_14 <= frequency_13;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_15 <= io_inputs_sortedFrequency_15;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_364) begin
            frequency_15 <= newFrequency;
          end else if (_T_365) begin
            frequency_15 <= frequency_14;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_16 <= io_inputs_sortedFrequency_16;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_366) begin
            frequency_16 <= newFrequency;
          end else if (_T_367) begin
            frequency_16 <= frequency_15;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_17 <= io_inputs_sortedFrequency_17;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_368) begin
            frequency_17 <= newFrequency;
          end else if (_T_369) begin
            frequency_17 <= frequency_16;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_18 <= io_inputs_sortedFrequency_18;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_370) begin
            frequency_18 <= newFrequency;
          end else if (_T_371) begin
            frequency_18 <= frequency_17;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_19 <= io_inputs_sortedFrequency_19;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_372) begin
            frequency_19 <= newFrequency;
          end else if (_T_373) begin
            frequency_19 <= frequency_18;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_20 <= io_inputs_sortedFrequency_20;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_374) begin
            frequency_20 <= newFrequency;
          end else if (_T_375) begin
            frequency_20 <= frequency_19;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_21 <= io_inputs_sortedFrequency_21;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_376) begin
            frequency_21 <= newFrequency;
          end else if (_T_377) begin
            frequency_21 <= frequency_20;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_22 <= io_inputs_sortedFrequency_22;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_378) begin
            frequency_22 <= newFrequency;
          end else if (_T_379) begin
            frequency_22 <= frequency_21;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_23 <= io_inputs_sortedFrequency_23;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_380) begin
            frequency_23 <= newFrequency;
          end else if (_T_381) begin
            frequency_23 <= frequency_22;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_24 <= io_inputs_sortedFrequency_24;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_382) begin
            frequency_24 <= newFrequency;
          end else if (_T_383) begin
            frequency_24 <= frequency_23;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_25 <= io_inputs_sortedFrequency_25;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_384) begin
            frequency_25 <= newFrequency;
          end else if (_T_385) begin
            frequency_25 <= frequency_24;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_26 <= io_inputs_sortedFrequency_26;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_386) begin
            frequency_26 <= newFrequency;
          end else if (_T_387) begin
            frequency_26 <= frequency_25;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_27 <= io_inputs_sortedFrequency_27;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_388) begin
            frequency_27 <= newFrequency;
          end else if (_T_389) begin
            frequency_27 <= frequency_26;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_28 <= io_inputs_sortedFrequency_28;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_390) begin
            frequency_28 <= newFrequency;
          end else if (_T_391) begin
            frequency_28 <= frequency_27;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_29 <= io_inputs_sortedFrequency_29;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_392) begin
            frequency_29 <= newFrequency;
          end else if (_T_393) begin
            frequency_29 <= frequency_28;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_30 <= io_inputs_sortedFrequency_30;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_394) begin
            frequency_30 <= newFrequency;
          end else if (_T_395) begin
            frequency_30 <= frequency_29;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        frequency_31 <= io_inputs_sortedFrequency_31;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_396) begin
            frequency_31 <= newFrequency;
          end else if (_T_397) begin
            frequency_31 <= frequency_30;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_0 <= io_inputs_sortedCharacter_0;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_334) begin
            pointerOrCharacter_0 <= newPointer;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_1 <= io_inputs_sortedCharacter_1;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_336) begin
            pointerOrCharacter_1 <= newPointer;
          end else if (_T_337) begin
            pointerOrCharacter_1 <= pointerOrCharacter_0;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_2 <= io_inputs_sortedCharacter_2;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_338) begin
            pointerOrCharacter_2 <= newPointer;
          end else if (_T_339) begin
            pointerOrCharacter_2 <= pointerOrCharacter_1;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_3 <= io_inputs_sortedCharacter_3;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_340) begin
            pointerOrCharacter_3 <= newPointer;
          end else if (_T_341) begin
            pointerOrCharacter_3 <= pointerOrCharacter_2;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_4 <= io_inputs_sortedCharacter_4;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_342) begin
            pointerOrCharacter_4 <= newPointer;
          end else if (_T_343) begin
            pointerOrCharacter_4 <= pointerOrCharacter_3;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_5 <= io_inputs_sortedCharacter_5;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_344) begin
            pointerOrCharacter_5 <= newPointer;
          end else if (_T_345) begin
            pointerOrCharacter_5 <= pointerOrCharacter_4;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_6 <= io_inputs_sortedCharacter_6;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_346) begin
            pointerOrCharacter_6 <= newPointer;
          end else if (_T_347) begin
            pointerOrCharacter_6 <= pointerOrCharacter_5;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_7 <= io_inputs_sortedCharacter_7;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_348) begin
            pointerOrCharacter_7 <= newPointer;
          end else if (_T_349) begin
            pointerOrCharacter_7 <= pointerOrCharacter_6;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_8 <= io_inputs_sortedCharacter_8;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_350) begin
            pointerOrCharacter_8 <= newPointer;
          end else if (_T_351) begin
            pointerOrCharacter_8 <= pointerOrCharacter_7;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_9 <= io_inputs_sortedCharacter_9;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_352) begin
            pointerOrCharacter_9 <= newPointer;
          end else if (_T_353) begin
            pointerOrCharacter_9 <= pointerOrCharacter_8;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_10 <= io_inputs_sortedCharacter_10;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_354) begin
            pointerOrCharacter_10 <= newPointer;
          end else if (_T_355) begin
            pointerOrCharacter_10 <= pointerOrCharacter_9;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_11 <= io_inputs_sortedCharacter_11;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_356) begin
            pointerOrCharacter_11 <= newPointer;
          end else if (_T_357) begin
            pointerOrCharacter_11 <= pointerOrCharacter_10;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_12 <= io_inputs_sortedCharacter_12;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_358) begin
            pointerOrCharacter_12 <= newPointer;
          end else if (_T_359) begin
            pointerOrCharacter_12 <= pointerOrCharacter_11;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_13 <= io_inputs_sortedCharacter_13;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_360) begin
            pointerOrCharacter_13 <= newPointer;
          end else if (_T_361) begin
            pointerOrCharacter_13 <= pointerOrCharacter_12;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_14 <= io_inputs_sortedCharacter_14;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_362) begin
            pointerOrCharacter_14 <= newPointer;
          end else if (_T_363) begin
            pointerOrCharacter_14 <= pointerOrCharacter_13;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_15 <= io_inputs_sortedCharacter_15;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_364) begin
            pointerOrCharacter_15 <= newPointer;
          end else if (_T_365) begin
            pointerOrCharacter_15 <= pointerOrCharacter_14;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_16 <= io_inputs_sortedCharacter_16;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_366) begin
            pointerOrCharacter_16 <= newPointer;
          end else if (_T_367) begin
            pointerOrCharacter_16 <= pointerOrCharacter_15;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_17 <= io_inputs_sortedCharacter_17;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_368) begin
            pointerOrCharacter_17 <= newPointer;
          end else if (_T_369) begin
            pointerOrCharacter_17 <= pointerOrCharacter_16;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_18 <= io_inputs_sortedCharacter_18;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_370) begin
            pointerOrCharacter_18 <= newPointer;
          end else if (_T_371) begin
            pointerOrCharacter_18 <= pointerOrCharacter_17;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_19 <= io_inputs_sortedCharacter_19;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_372) begin
            pointerOrCharacter_19 <= newPointer;
          end else if (_T_373) begin
            pointerOrCharacter_19 <= pointerOrCharacter_18;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_20 <= io_inputs_sortedCharacter_20;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_374) begin
            pointerOrCharacter_20 <= newPointer;
          end else if (_T_375) begin
            pointerOrCharacter_20 <= pointerOrCharacter_19;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_21 <= io_inputs_sortedCharacter_21;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_376) begin
            pointerOrCharacter_21 <= newPointer;
          end else if (_T_377) begin
            pointerOrCharacter_21 <= pointerOrCharacter_20;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_22 <= io_inputs_sortedCharacter_22;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_378) begin
            pointerOrCharacter_22 <= newPointer;
          end else if (_T_379) begin
            pointerOrCharacter_22 <= pointerOrCharacter_21;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_23 <= io_inputs_sortedCharacter_23;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_380) begin
            pointerOrCharacter_23 <= newPointer;
          end else if (_T_381) begin
            pointerOrCharacter_23 <= pointerOrCharacter_22;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_24 <= io_inputs_sortedCharacter_24;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_382) begin
            pointerOrCharacter_24 <= newPointer;
          end else if (_T_383) begin
            pointerOrCharacter_24 <= pointerOrCharacter_23;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_25 <= io_inputs_sortedCharacter_25;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_384) begin
            pointerOrCharacter_25 <= newPointer;
          end else if (_T_385) begin
            pointerOrCharacter_25 <= pointerOrCharacter_24;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_26 <= io_inputs_sortedCharacter_26;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_386) begin
            pointerOrCharacter_26 <= newPointer;
          end else if (_T_387) begin
            pointerOrCharacter_26 <= pointerOrCharacter_25;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_27 <= io_inputs_sortedCharacter_27;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_388) begin
            pointerOrCharacter_27 <= newPointer;
          end else if (_T_389) begin
            pointerOrCharacter_27 <= pointerOrCharacter_26;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_28 <= io_inputs_sortedCharacter_28;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_390) begin
            pointerOrCharacter_28 <= newPointer;
          end else if (_T_391) begin
            pointerOrCharacter_28 <= pointerOrCharacter_27;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_29 <= io_inputs_sortedCharacter_29;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_392) begin
            pointerOrCharacter_29 <= newPointer;
          end else if (_T_393) begin
            pointerOrCharacter_29 <= pointerOrCharacter_28;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_30 <= io_inputs_sortedCharacter_30;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_394) begin
            pointerOrCharacter_30 <= newPointer;
          end else if (_T_395) begin
            pointerOrCharacter_30 <= pointerOrCharacter_29;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        pointerOrCharacter_31 <= io_inputs_sortedCharacter_31;
      end
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_396) begin
            pointerOrCharacter_31 <= newPointer;
          end else if (_T_397) begin
            pointerOrCharacter_31 <= pointerOrCharacter_30;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_0 <= _GEN_66;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_334) begin
            isCharacter_0 <= 1'h0;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_1 <= _GEN_67;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_336) begin
            isCharacter_1 <= 1'h0;
          end else if (_T_337) begin
            isCharacter_1 <= isCharacter_0;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_2 <= _GEN_68;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_338) begin
            isCharacter_2 <= 1'h0;
          end else if (_T_339) begin
            isCharacter_2 <= isCharacter_1;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_3 <= _GEN_69;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_340) begin
            isCharacter_3 <= 1'h0;
          end else if (_T_341) begin
            isCharacter_3 <= isCharacter_2;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_4 <= _GEN_70;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_342) begin
            isCharacter_4 <= 1'h0;
          end else if (_T_343) begin
            isCharacter_4 <= isCharacter_3;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_5 <= _GEN_71;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_344) begin
            isCharacter_5 <= 1'h0;
          end else if (_T_345) begin
            isCharacter_5 <= isCharacter_4;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_6 <= _GEN_72;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_346) begin
            isCharacter_6 <= 1'h0;
          end else if (_T_347) begin
            isCharacter_6 <= isCharacter_5;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_7 <= _GEN_73;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_348) begin
            isCharacter_7 <= 1'h0;
          end else if (_T_349) begin
            isCharacter_7 <= isCharacter_6;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_8 <= _GEN_74;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_350) begin
            isCharacter_8 <= 1'h0;
          end else if (_T_351) begin
            isCharacter_8 <= isCharacter_7;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_9 <= _GEN_75;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_352) begin
            isCharacter_9 <= 1'h0;
          end else if (_T_353) begin
            isCharacter_9 <= isCharacter_8;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_10 <= _GEN_76;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_354) begin
            isCharacter_10 <= 1'h0;
          end else if (_T_355) begin
            isCharacter_10 <= isCharacter_9;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_11 <= _GEN_77;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_356) begin
            isCharacter_11 <= 1'h0;
          end else if (_T_357) begin
            isCharacter_11 <= isCharacter_10;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_12 <= _GEN_78;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_358) begin
            isCharacter_12 <= 1'h0;
          end else if (_T_359) begin
            isCharacter_12 <= isCharacter_11;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_13 <= _GEN_79;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_360) begin
            isCharacter_13 <= 1'h0;
          end else if (_T_361) begin
            isCharacter_13 <= isCharacter_12;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_14 <= _GEN_80;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_362) begin
            isCharacter_14 <= 1'h0;
          end else if (_T_363) begin
            isCharacter_14 <= isCharacter_13;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_15 <= _GEN_81;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_364) begin
            isCharacter_15 <= 1'h0;
          end else if (_T_365) begin
            isCharacter_15 <= isCharacter_14;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_16 <= _GEN_82;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_366) begin
            isCharacter_16 <= 1'h0;
          end else if (_T_367) begin
            isCharacter_16 <= isCharacter_15;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_17 <= _GEN_83;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_368) begin
            isCharacter_17 <= 1'h0;
          end else if (_T_369) begin
            isCharacter_17 <= isCharacter_16;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_18 <= _GEN_84;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_370) begin
            isCharacter_18 <= 1'h0;
          end else if (_T_371) begin
            isCharacter_18 <= isCharacter_17;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_19 <= _GEN_85;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_372) begin
            isCharacter_19 <= 1'h0;
          end else if (_T_373) begin
            isCharacter_19 <= isCharacter_18;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_20 <= _GEN_86;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_374) begin
            isCharacter_20 <= 1'h0;
          end else if (_T_375) begin
            isCharacter_20 <= isCharacter_19;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_21 <= _GEN_87;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_376) begin
            isCharacter_21 <= 1'h0;
          end else if (_T_377) begin
            isCharacter_21 <= isCharacter_20;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_22 <= _GEN_88;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_378) begin
            isCharacter_22 <= 1'h0;
          end else if (_T_379) begin
            isCharacter_22 <= isCharacter_21;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_23 <= _GEN_89;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_380) begin
            isCharacter_23 <= 1'h0;
          end else if (_T_381) begin
            isCharacter_23 <= isCharacter_22;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_24 <= _GEN_90;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_382) begin
            isCharacter_24 <= 1'h0;
          end else if (_T_383) begin
            isCharacter_24 <= isCharacter_23;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_25 <= _GEN_91;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_384) begin
            isCharacter_25 <= 1'h0;
          end else if (_T_385) begin
            isCharacter_25 <= isCharacter_24;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_26 <= _GEN_92;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_386) begin
            isCharacter_26 <= 1'h0;
          end else if (_T_387) begin
            isCharacter_26 <= isCharacter_25;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_27 <= _GEN_93;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_388) begin
            isCharacter_27 <= 1'h0;
          end else if (_T_389) begin
            isCharacter_27 <= isCharacter_26;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_28 <= _GEN_94;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_390) begin
            isCharacter_28 <= 1'h0;
          end else if (_T_391) begin
            isCharacter_28 <= isCharacter_27;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_29 <= _GEN_95;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_392) begin
            isCharacter_29 <= 1'h0;
          end else if (_T_393) begin
            isCharacter_29 <= isCharacter_28;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_30 <= _GEN_96;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_394) begin
            isCharacter_30 <= 1'h0;
          end else if (_T_395) begin
            isCharacter_30 <= isCharacter_29;
          end
        end
      end
    end
    if (_T_32) begin
      isCharacter_31 <= _GEN_97;
    end else if (!(_T_284)) begin
      if (_T_317) begin
        if (searchCompleted) begin
          if (_T_396) begin
            isCharacter_31 <= 1'h0;
          end else if (_T_397) begin
            isCharacter_31 <= isCharacter_30;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          newFrequency <= _T_314;
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          newPointer <= {{2'd0}, validNodes};
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        validRoots <= _T_157;
      end
    end else if (_T_284) begin
      if (!(_T_285)) begin
        validRoots <= _T_290;
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (_T_285) begin
          if (_T_286) begin
            leftNode_0 <= pointerOrCharacter_0;
          end
        end else if (6'h0 == validNodes[5:0]) begin
          if (5'h1f == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_31;
          end else if (5'h1e == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_30;
          end else if (5'h1d == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_29;
          end else if (5'h1c == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_28;
          end else if (5'h1b == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_27;
          end else if (5'h1a == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_26;
          end else if (5'h19 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_25;
          end else if (5'h18 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_24;
          end else if (5'h17 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_23;
          end else if (5'h16 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_22;
          end else if (5'h15 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_21;
          end else if (5'h14 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_20;
          end else if (5'h13 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_19;
          end else if (5'h12 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_18;
          end else if (5'h11 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_17;
          end else if (5'h10 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_16;
          end else if (5'hf == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_15;
          end else if (5'he == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_14;
          end else if (5'hd == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_13;
          end else if (5'hc == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_12;
          end else if (5'hb == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_11;
          end else if (5'ha == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_10;
          end else if (5'h9 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_9;
          end else if (5'h8 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_8;
          end else if (5'h7 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_7;
          end else if (5'h6 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_6;
          end else if (5'h5 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_5;
          end else if (5'h4 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_4;
          end else if (5'h3 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_3;
          end else if (5'h2 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_2;
          end else if (5'h1 == _T_293[4:0]) begin
            leftNode_0 <= pointerOrCharacter_1;
          end else begin
            leftNode_0 <= pointerOrCharacter_0;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1 == validNodes[5:0]) begin
            if (5'h1f == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_31;
            end else if (5'h1e == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_30;
            end else if (5'h1d == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_29;
            end else if (5'h1c == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_28;
            end else if (5'h1b == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_27;
            end else if (5'h1a == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_26;
            end else if (5'h19 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_25;
            end else if (5'h18 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_24;
            end else if (5'h17 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_23;
            end else if (5'h16 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_22;
            end else if (5'h15 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_21;
            end else if (5'h14 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_20;
            end else if (5'h13 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_19;
            end else if (5'h12 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_18;
            end else if (5'h11 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_17;
            end else if (5'h10 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_16;
            end else if (5'hf == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_15;
            end else if (5'he == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_14;
            end else if (5'hd == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_13;
            end else if (5'hc == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_12;
            end else if (5'hb == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_11;
            end else if (5'ha == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_10;
            end else if (5'h9 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_9;
            end else if (5'h8 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_8;
            end else if (5'h7 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_7;
            end else if (5'h6 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_6;
            end else if (5'h5 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_5;
            end else if (5'h4 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_4;
            end else if (5'h3 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_3;
            end else if (5'h2 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_2;
            end else if (5'h1 == _T_293[4:0]) begin
              leftNode_1 <= pointerOrCharacter_1;
            end else begin
              leftNode_1 <= pointerOrCharacter_0;
            end
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2 == validNodes[5:0]) begin
            if (5'h1f == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_31;
            end else if (5'h1e == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_30;
            end else if (5'h1d == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_29;
            end else if (5'h1c == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_28;
            end else if (5'h1b == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_27;
            end else if (5'h1a == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_26;
            end else if (5'h19 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_25;
            end else if (5'h18 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_24;
            end else if (5'h17 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_23;
            end else if (5'h16 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_22;
            end else if (5'h15 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_21;
            end else if (5'h14 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_20;
            end else if (5'h13 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_19;
            end else if (5'h12 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_18;
            end else if (5'h11 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_17;
            end else if (5'h10 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_16;
            end else if (5'hf == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_15;
            end else if (5'he == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_14;
            end else if (5'hd == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_13;
            end else if (5'hc == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_12;
            end else if (5'hb == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_11;
            end else if (5'ha == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_10;
            end else if (5'h9 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_9;
            end else if (5'h8 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_8;
            end else if (5'h7 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_7;
            end else if (5'h6 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_6;
            end else if (5'h5 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_5;
            end else if (5'h4 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_4;
            end else if (5'h3 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_3;
            end else if (5'h2 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_2;
            end else if (5'h1 == _T_293[4:0]) begin
              leftNode_2 <= pointerOrCharacter_1;
            end else begin
              leftNode_2 <= pointerOrCharacter_0;
            end
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3 == validNodes[5:0]) begin
            if (5'h1f == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_31;
            end else if (5'h1e == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_30;
            end else if (5'h1d == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_29;
            end else if (5'h1c == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_28;
            end else if (5'h1b == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_27;
            end else if (5'h1a == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_26;
            end else if (5'h19 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_25;
            end else if (5'h18 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_24;
            end else if (5'h17 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_23;
            end else if (5'h16 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_22;
            end else if (5'h15 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_21;
            end else if (5'h14 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_20;
            end else if (5'h13 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_19;
            end else if (5'h12 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_18;
            end else if (5'h11 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_17;
            end else if (5'h10 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_16;
            end else if (5'hf == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_15;
            end else if (5'he == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_14;
            end else if (5'hd == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_13;
            end else if (5'hc == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_12;
            end else if (5'hb == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_11;
            end else if (5'ha == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_10;
            end else if (5'h9 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_9;
            end else if (5'h8 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_8;
            end else if (5'h7 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_7;
            end else if (5'h6 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_6;
            end else if (5'h5 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_5;
            end else if (5'h4 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_4;
            end else if (5'h3 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_3;
            end else if (5'h2 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_2;
            end else if (5'h1 == _T_293[4:0]) begin
              leftNode_3 <= pointerOrCharacter_1;
            end else begin
              leftNode_3 <= pointerOrCharacter_0;
            end
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h4 == validNodes[5:0]) begin
            leftNode_4 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h5 == validNodes[5:0]) begin
            leftNode_5 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h6 == validNodes[5:0]) begin
            leftNode_6 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h7 == validNodes[5:0]) begin
            leftNode_7 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h8 == validNodes[5:0]) begin
            leftNode_8 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h9 == validNodes[5:0]) begin
            leftNode_9 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'ha == validNodes[5:0]) begin
            leftNode_10 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'hb == validNodes[5:0]) begin
            leftNode_11 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'hc == validNodes[5:0]) begin
            leftNode_12 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'hd == validNodes[5:0]) begin
            leftNode_13 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'he == validNodes[5:0]) begin
            leftNode_14 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'hf == validNodes[5:0]) begin
            leftNode_15 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h10 == validNodes[5:0]) begin
            leftNode_16 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h11 == validNodes[5:0]) begin
            leftNode_17 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h12 == validNodes[5:0]) begin
            leftNode_18 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h13 == validNodes[5:0]) begin
            leftNode_19 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h14 == validNodes[5:0]) begin
            leftNode_20 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h15 == validNodes[5:0]) begin
            leftNode_21 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h16 == validNodes[5:0]) begin
            leftNode_22 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h17 == validNodes[5:0]) begin
            leftNode_23 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h18 == validNodes[5:0]) begin
            leftNode_24 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h19 == validNodes[5:0]) begin
            leftNode_25 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1a == validNodes[5:0]) begin
            leftNode_26 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1b == validNodes[5:0]) begin
            leftNode_27 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1c == validNodes[5:0]) begin
            leftNode_28 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1d == validNodes[5:0]) begin
            leftNode_29 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1e == validNodes[5:0]) begin
            leftNode_30 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1f == validNodes[5:0]) begin
            leftNode_31 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h20 == validNodes[5:0]) begin
            leftNode_32 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h21 == validNodes[5:0]) begin
            leftNode_33 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h22 == validNodes[5:0]) begin
            leftNode_34 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h23 == validNodes[5:0]) begin
            leftNode_35 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h24 == validNodes[5:0]) begin
            leftNode_36 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h25 == validNodes[5:0]) begin
            leftNode_37 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h26 == validNodes[5:0]) begin
            leftNode_38 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h27 == validNodes[5:0]) begin
            leftNode_39 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h28 == validNodes[5:0]) begin
            leftNode_40 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h29 == validNodes[5:0]) begin
            leftNode_41 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2a == validNodes[5:0]) begin
            leftNode_42 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2b == validNodes[5:0]) begin
            leftNode_43 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2c == validNodes[5:0]) begin
            leftNode_44 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2d == validNodes[5:0]) begin
            leftNode_45 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2e == validNodes[5:0]) begin
            leftNode_46 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2f == validNodes[5:0]) begin
            leftNode_47 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h30 == validNodes[5:0]) begin
            leftNode_48 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h31 == validNodes[5:0]) begin
            leftNode_49 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h32 == validNodes[5:0]) begin
            leftNode_50 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h33 == validNodes[5:0]) begin
            leftNode_51 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h34 == validNodes[5:0]) begin
            leftNode_52 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h35 == validNodes[5:0]) begin
            leftNode_53 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h36 == validNodes[5:0]) begin
            leftNode_54 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h37 == validNodes[5:0]) begin
            leftNode_55 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h38 == validNodes[5:0]) begin
            leftNode_56 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h39 == validNodes[5:0]) begin
            leftNode_57 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3a == validNodes[5:0]) begin
            leftNode_58 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3b == validNodes[5:0]) begin
            leftNode_59 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3c == validNodes[5:0]) begin
            leftNode_60 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3d == validNodes[5:0]) begin
            leftNode_61 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3e == validNodes[5:0]) begin
            leftNode_62 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3f == validNodes[5:0]) begin
            leftNode_63 <= _GEN_199;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h0 == validNodes[5:0]) begin
            if (5'h1f == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_31;
            end else if (5'h1e == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_30;
            end else if (5'h1d == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_29;
            end else if (5'h1c == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_28;
            end else if (5'h1b == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_27;
            end else if (5'h1a == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_26;
            end else if (5'h19 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_25;
            end else if (5'h18 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_24;
            end else if (5'h17 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_23;
            end else if (5'h16 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_22;
            end else if (5'h15 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_21;
            end else if (5'h14 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_20;
            end else if (5'h13 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_19;
            end else if (5'h12 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_18;
            end else if (5'h11 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_17;
            end else if (5'h10 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_16;
            end else if (5'hf == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_15;
            end else if (5'he == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_14;
            end else if (5'hd == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_13;
            end else if (5'hc == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_12;
            end else if (5'hb == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_11;
            end else if (5'ha == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_10;
            end else if (5'h9 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_9;
            end else if (5'h8 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_8;
            end else if (5'h7 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_7;
            end else if (5'h6 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_6;
            end else if (5'h5 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_5;
            end else if (5'h4 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_4;
            end else if (5'h3 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_3;
            end else if (5'h2 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_2;
            end else if (5'h1 == _T_290[4:0]) begin
              rightNode_0 <= pointerOrCharacter_1;
            end else begin
              rightNode_0 <= pointerOrCharacter_0;
            end
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1 == validNodes[5:0]) begin
            if (5'h1f == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_31;
            end else if (5'h1e == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_30;
            end else if (5'h1d == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_29;
            end else if (5'h1c == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_28;
            end else if (5'h1b == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_27;
            end else if (5'h1a == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_26;
            end else if (5'h19 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_25;
            end else if (5'h18 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_24;
            end else if (5'h17 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_23;
            end else if (5'h16 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_22;
            end else if (5'h15 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_21;
            end else if (5'h14 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_20;
            end else if (5'h13 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_19;
            end else if (5'h12 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_18;
            end else if (5'h11 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_17;
            end else if (5'h10 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_16;
            end else if (5'hf == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_15;
            end else if (5'he == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_14;
            end else if (5'hd == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_13;
            end else if (5'hc == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_12;
            end else if (5'hb == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_11;
            end else if (5'ha == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_10;
            end else if (5'h9 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_9;
            end else if (5'h8 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_8;
            end else if (5'h7 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_7;
            end else if (5'h6 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_6;
            end else if (5'h5 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_5;
            end else if (5'h4 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_4;
            end else if (5'h3 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_3;
            end else if (5'h2 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_2;
            end else if (5'h1 == _T_290[4:0]) begin
              rightNode_1 <= pointerOrCharacter_1;
            end else begin
              rightNode_1 <= pointerOrCharacter_0;
            end
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2 == validNodes[5:0]) begin
            if (5'h1f == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_31;
            end else if (5'h1e == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_30;
            end else if (5'h1d == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_29;
            end else if (5'h1c == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_28;
            end else if (5'h1b == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_27;
            end else if (5'h1a == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_26;
            end else if (5'h19 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_25;
            end else if (5'h18 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_24;
            end else if (5'h17 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_23;
            end else if (5'h16 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_22;
            end else if (5'h15 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_21;
            end else if (5'h14 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_20;
            end else if (5'h13 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_19;
            end else if (5'h12 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_18;
            end else if (5'h11 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_17;
            end else if (5'h10 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_16;
            end else if (5'hf == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_15;
            end else if (5'he == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_14;
            end else if (5'hd == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_13;
            end else if (5'hc == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_12;
            end else if (5'hb == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_11;
            end else if (5'ha == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_10;
            end else if (5'h9 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_9;
            end else if (5'h8 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_8;
            end else if (5'h7 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_7;
            end else if (5'h6 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_6;
            end else if (5'h5 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_5;
            end else if (5'h4 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_4;
            end else if (5'h3 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_3;
            end else if (5'h2 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_2;
            end else if (5'h1 == _T_290[4:0]) begin
              rightNode_2 <= pointerOrCharacter_1;
            end else begin
              rightNode_2 <= pointerOrCharacter_0;
            end
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3 == validNodes[5:0]) begin
            if (5'h1f == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_31;
            end else if (5'h1e == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_30;
            end else if (5'h1d == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_29;
            end else if (5'h1c == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_28;
            end else if (5'h1b == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_27;
            end else if (5'h1a == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_26;
            end else if (5'h19 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_25;
            end else if (5'h18 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_24;
            end else if (5'h17 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_23;
            end else if (5'h16 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_22;
            end else if (5'h15 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_21;
            end else if (5'h14 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_20;
            end else if (5'h13 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_19;
            end else if (5'h12 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_18;
            end else if (5'h11 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_17;
            end else if (5'h10 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_16;
            end else if (5'hf == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_15;
            end else if (5'he == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_14;
            end else if (5'hd == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_13;
            end else if (5'hc == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_12;
            end else if (5'hb == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_11;
            end else if (5'ha == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_10;
            end else if (5'h9 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_9;
            end else if (5'h8 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_8;
            end else if (5'h7 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_7;
            end else if (5'h6 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_6;
            end else if (5'h5 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_5;
            end else if (5'h4 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_4;
            end else if (5'h3 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_3;
            end else if (5'h2 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_2;
            end else if (5'h1 == _T_290[4:0]) begin
              rightNode_3 <= pointerOrCharacter_1;
            end else begin
              rightNode_3 <= pointerOrCharacter_0;
            end
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h4 == validNodes[5:0]) begin
            rightNode_4 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h5 == validNodes[5:0]) begin
            rightNode_5 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h6 == validNodes[5:0]) begin
            rightNode_6 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h7 == validNodes[5:0]) begin
            rightNode_7 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h8 == validNodes[5:0]) begin
            rightNode_8 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h9 == validNodes[5:0]) begin
            rightNode_9 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'ha == validNodes[5:0]) begin
            rightNode_10 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'hb == validNodes[5:0]) begin
            rightNode_11 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'hc == validNodes[5:0]) begin
            rightNode_12 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'hd == validNodes[5:0]) begin
            rightNode_13 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'he == validNodes[5:0]) begin
            rightNode_14 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'hf == validNodes[5:0]) begin
            rightNode_15 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h10 == validNodes[5:0]) begin
            rightNode_16 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h11 == validNodes[5:0]) begin
            rightNode_17 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h12 == validNodes[5:0]) begin
            rightNode_18 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h13 == validNodes[5:0]) begin
            rightNode_19 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h14 == validNodes[5:0]) begin
            rightNode_20 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h15 == validNodes[5:0]) begin
            rightNode_21 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h16 == validNodes[5:0]) begin
            rightNode_22 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h17 == validNodes[5:0]) begin
            rightNode_23 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h18 == validNodes[5:0]) begin
            rightNode_24 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h19 == validNodes[5:0]) begin
            rightNode_25 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1a == validNodes[5:0]) begin
            rightNode_26 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1b == validNodes[5:0]) begin
            rightNode_27 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1c == validNodes[5:0]) begin
            rightNode_28 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1d == validNodes[5:0]) begin
            rightNode_29 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1e == validNodes[5:0]) begin
            rightNode_30 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1f == validNodes[5:0]) begin
            rightNode_31 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h20 == validNodes[5:0]) begin
            rightNode_32 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h21 == validNodes[5:0]) begin
            rightNode_33 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h22 == validNodes[5:0]) begin
            rightNode_34 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h23 == validNodes[5:0]) begin
            rightNode_35 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h24 == validNodes[5:0]) begin
            rightNode_36 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h25 == validNodes[5:0]) begin
            rightNode_37 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h26 == validNodes[5:0]) begin
            rightNode_38 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h27 == validNodes[5:0]) begin
            rightNode_39 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h28 == validNodes[5:0]) begin
            rightNode_40 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h29 == validNodes[5:0]) begin
            rightNode_41 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2a == validNodes[5:0]) begin
            rightNode_42 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2b == validNodes[5:0]) begin
            rightNode_43 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2c == validNodes[5:0]) begin
            rightNode_44 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2d == validNodes[5:0]) begin
            rightNode_45 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2e == validNodes[5:0]) begin
            rightNode_46 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2f == validNodes[5:0]) begin
            rightNode_47 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h30 == validNodes[5:0]) begin
            rightNode_48 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h31 == validNodes[5:0]) begin
            rightNode_49 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h32 == validNodes[5:0]) begin
            rightNode_50 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h33 == validNodes[5:0]) begin
            rightNode_51 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h34 == validNodes[5:0]) begin
            rightNode_52 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h35 == validNodes[5:0]) begin
            rightNode_53 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h36 == validNodes[5:0]) begin
            rightNode_54 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h37 == validNodes[5:0]) begin
            rightNode_55 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h38 == validNodes[5:0]) begin
            rightNode_56 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h39 == validNodes[5:0]) begin
            rightNode_57 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3a == validNodes[5:0]) begin
            rightNode_58 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3b == validNodes[5:0]) begin
            rightNode_59 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3c == validNodes[5:0]) begin
            rightNode_60 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3d == validNodes[5:0]) begin
            rightNode_61 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3e == validNodes[5:0]) begin
            rightNode_62 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3f == validNodes[5:0]) begin
            rightNode_63 <= _GEN_391;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (_T_285) begin
          leftNodeIsCharacter_0 <= _GEN_103;
        end else if (6'h0 == validNodes[5:0]) begin
          if (5'h1f == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_31;
          end else if (5'h1e == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_30;
          end else if (5'h1d == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_29;
          end else if (5'h1c == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_28;
          end else if (5'h1b == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_27;
          end else if (5'h1a == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_26;
          end else if (5'h19 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_25;
          end else if (5'h18 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_24;
          end else if (5'h17 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_23;
          end else if (5'h16 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_22;
          end else if (5'h15 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_21;
          end else if (5'h14 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_20;
          end else if (5'h13 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_19;
          end else if (5'h12 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_18;
          end else if (5'h11 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_17;
          end else if (5'h10 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_16;
          end else if (5'hf == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_15;
          end else if (5'he == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_14;
          end else if (5'hd == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_13;
          end else if (5'hc == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_12;
          end else if (5'hb == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_11;
          end else if (5'ha == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_10;
          end else if (5'h9 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_9;
          end else if (5'h8 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_8;
          end else if (5'h7 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_7;
          end else if (5'h6 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_6;
          end else if (5'h5 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_5;
          end else if (5'h4 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_4;
          end else if (5'h3 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_3;
          end else if (5'h2 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_2;
          end else if (5'h1 == _T_293[4:0]) begin
            leftNodeIsCharacter_0 <= isCharacter_1;
          end else begin
            leftNodeIsCharacter_0 <= isCharacter_0;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1 == validNodes[5:0]) begin
            if (5'h1f == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_31;
            end else if (5'h1e == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_30;
            end else if (5'h1d == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_29;
            end else if (5'h1c == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_28;
            end else if (5'h1b == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_27;
            end else if (5'h1a == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_26;
            end else if (5'h19 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_25;
            end else if (5'h18 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_24;
            end else if (5'h17 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_23;
            end else if (5'h16 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_22;
            end else if (5'h15 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_21;
            end else if (5'h14 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_20;
            end else if (5'h13 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_19;
            end else if (5'h12 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_18;
            end else if (5'h11 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_17;
            end else if (5'h10 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_16;
            end else if (5'hf == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_15;
            end else if (5'he == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_14;
            end else if (5'hd == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_13;
            end else if (5'hc == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_12;
            end else if (5'hb == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_11;
            end else if (5'ha == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_10;
            end else if (5'h9 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_9;
            end else if (5'h8 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_8;
            end else if (5'h7 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_7;
            end else if (5'h6 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_6;
            end else if (5'h5 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_5;
            end else if (5'h4 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_4;
            end else if (5'h3 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_3;
            end else if (5'h2 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_2;
            end else if (5'h1 == _T_293[4:0]) begin
              leftNodeIsCharacter_1 <= isCharacter_1;
            end else begin
              leftNodeIsCharacter_1 <= isCharacter_0;
            end
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2 == validNodes[5:0]) begin
            if (5'h1f == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_31;
            end else if (5'h1e == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_30;
            end else if (5'h1d == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_29;
            end else if (5'h1c == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_28;
            end else if (5'h1b == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_27;
            end else if (5'h1a == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_26;
            end else if (5'h19 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_25;
            end else if (5'h18 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_24;
            end else if (5'h17 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_23;
            end else if (5'h16 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_22;
            end else if (5'h15 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_21;
            end else if (5'h14 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_20;
            end else if (5'h13 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_19;
            end else if (5'h12 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_18;
            end else if (5'h11 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_17;
            end else if (5'h10 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_16;
            end else if (5'hf == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_15;
            end else if (5'he == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_14;
            end else if (5'hd == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_13;
            end else if (5'hc == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_12;
            end else if (5'hb == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_11;
            end else if (5'ha == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_10;
            end else if (5'h9 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_9;
            end else if (5'h8 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_8;
            end else if (5'h7 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_7;
            end else if (5'h6 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_6;
            end else if (5'h5 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_5;
            end else if (5'h4 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_4;
            end else if (5'h3 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_3;
            end else if (5'h2 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_2;
            end else if (5'h1 == _T_293[4:0]) begin
              leftNodeIsCharacter_2 <= isCharacter_1;
            end else begin
              leftNodeIsCharacter_2 <= isCharacter_0;
            end
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3 == validNodes[5:0]) begin
            if (5'h1f == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_31;
            end else if (5'h1e == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_30;
            end else if (5'h1d == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_29;
            end else if (5'h1c == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_28;
            end else if (5'h1b == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_27;
            end else if (5'h1a == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_26;
            end else if (5'h19 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_25;
            end else if (5'h18 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_24;
            end else if (5'h17 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_23;
            end else if (5'h16 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_22;
            end else if (5'h15 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_21;
            end else if (5'h14 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_20;
            end else if (5'h13 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_19;
            end else if (5'h12 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_18;
            end else if (5'h11 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_17;
            end else if (5'h10 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_16;
            end else if (5'hf == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_15;
            end else if (5'he == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_14;
            end else if (5'hd == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_13;
            end else if (5'hc == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_12;
            end else if (5'hb == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_11;
            end else if (5'ha == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_10;
            end else if (5'h9 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_9;
            end else if (5'h8 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_8;
            end else if (5'h7 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_7;
            end else if (5'h6 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_6;
            end else if (5'h5 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_5;
            end else if (5'h4 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_4;
            end else if (5'h3 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_3;
            end else if (5'h2 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_2;
            end else if (5'h1 == _T_293[4:0]) begin
              leftNodeIsCharacter_3 <= isCharacter_1;
            end else begin
              leftNodeIsCharacter_3 <= isCharacter_0;
            end
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h4 == validNodes[5:0]) begin
            leftNodeIsCharacter_4 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h5 == validNodes[5:0]) begin
            leftNodeIsCharacter_5 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h6 == validNodes[5:0]) begin
            leftNodeIsCharacter_6 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h7 == validNodes[5:0]) begin
            leftNodeIsCharacter_7 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h8 == validNodes[5:0]) begin
            leftNodeIsCharacter_8 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h9 == validNodes[5:0]) begin
            leftNodeIsCharacter_9 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'ha == validNodes[5:0]) begin
            leftNodeIsCharacter_10 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'hb == validNodes[5:0]) begin
            leftNodeIsCharacter_11 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'hc == validNodes[5:0]) begin
            leftNodeIsCharacter_12 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'hd == validNodes[5:0]) begin
            leftNodeIsCharacter_13 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'he == validNodes[5:0]) begin
            leftNodeIsCharacter_14 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'hf == validNodes[5:0]) begin
            leftNodeIsCharacter_15 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h10 == validNodes[5:0]) begin
            leftNodeIsCharacter_16 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h11 == validNodes[5:0]) begin
            leftNodeIsCharacter_17 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h12 == validNodes[5:0]) begin
            leftNodeIsCharacter_18 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h13 == validNodes[5:0]) begin
            leftNodeIsCharacter_19 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h14 == validNodes[5:0]) begin
            leftNodeIsCharacter_20 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h15 == validNodes[5:0]) begin
            leftNodeIsCharacter_21 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h16 == validNodes[5:0]) begin
            leftNodeIsCharacter_22 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h17 == validNodes[5:0]) begin
            leftNodeIsCharacter_23 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h18 == validNodes[5:0]) begin
            leftNodeIsCharacter_24 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h19 == validNodes[5:0]) begin
            leftNodeIsCharacter_25 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1a == validNodes[5:0]) begin
            leftNodeIsCharacter_26 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1b == validNodes[5:0]) begin
            leftNodeIsCharacter_27 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1c == validNodes[5:0]) begin
            leftNodeIsCharacter_28 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1d == validNodes[5:0]) begin
            leftNodeIsCharacter_29 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1e == validNodes[5:0]) begin
            leftNodeIsCharacter_30 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1f == validNodes[5:0]) begin
            leftNodeIsCharacter_31 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h20 == validNodes[5:0]) begin
            leftNodeIsCharacter_32 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h21 == validNodes[5:0]) begin
            leftNodeIsCharacter_33 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h22 == validNodes[5:0]) begin
            leftNodeIsCharacter_34 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h23 == validNodes[5:0]) begin
            leftNodeIsCharacter_35 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h24 == validNodes[5:0]) begin
            leftNodeIsCharacter_36 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h25 == validNodes[5:0]) begin
            leftNodeIsCharacter_37 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h26 == validNodes[5:0]) begin
            leftNodeIsCharacter_38 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h27 == validNodes[5:0]) begin
            leftNodeIsCharacter_39 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h28 == validNodes[5:0]) begin
            leftNodeIsCharacter_40 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h29 == validNodes[5:0]) begin
            leftNodeIsCharacter_41 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2a == validNodes[5:0]) begin
            leftNodeIsCharacter_42 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2b == validNodes[5:0]) begin
            leftNodeIsCharacter_43 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2c == validNodes[5:0]) begin
            leftNodeIsCharacter_44 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2d == validNodes[5:0]) begin
            leftNodeIsCharacter_45 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2e == validNodes[5:0]) begin
            leftNodeIsCharacter_46 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2f == validNodes[5:0]) begin
            leftNodeIsCharacter_47 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h30 == validNodes[5:0]) begin
            leftNodeIsCharacter_48 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h31 == validNodes[5:0]) begin
            leftNodeIsCharacter_49 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h32 == validNodes[5:0]) begin
            leftNodeIsCharacter_50 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h33 == validNodes[5:0]) begin
            leftNodeIsCharacter_51 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h34 == validNodes[5:0]) begin
            leftNodeIsCharacter_52 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h35 == validNodes[5:0]) begin
            leftNodeIsCharacter_53 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h36 == validNodes[5:0]) begin
            leftNodeIsCharacter_54 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h37 == validNodes[5:0]) begin
            leftNodeIsCharacter_55 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h38 == validNodes[5:0]) begin
            leftNodeIsCharacter_56 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h39 == validNodes[5:0]) begin
            leftNodeIsCharacter_57 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3a == validNodes[5:0]) begin
            leftNodeIsCharacter_58 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3b == validNodes[5:0]) begin
            leftNodeIsCharacter_59 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3c == validNodes[5:0]) begin
            leftNodeIsCharacter_60 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3d == validNodes[5:0]) begin
            leftNodeIsCharacter_61 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3e == validNodes[5:0]) begin
            leftNodeIsCharacter_62 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3f == validNodes[5:0]) begin
            leftNodeIsCharacter_63 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h0 == validNodes[5:0]) begin
            if (5'h1f == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_31;
            end else if (5'h1e == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_30;
            end else if (5'h1d == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_29;
            end else if (5'h1c == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_28;
            end else if (5'h1b == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_27;
            end else if (5'h1a == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_26;
            end else if (5'h19 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_25;
            end else if (5'h18 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_24;
            end else if (5'h17 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_23;
            end else if (5'h16 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_22;
            end else if (5'h15 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_21;
            end else if (5'h14 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_20;
            end else if (5'h13 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_19;
            end else if (5'h12 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_18;
            end else if (5'h11 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_17;
            end else if (5'h10 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_16;
            end else if (5'hf == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_15;
            end else if (5'he == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_14;
            end else if (5'hd == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_13;
            end else if (5'hc == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_12;
            end else if (5'hb == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_11;
            end else if (5'ha == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_10;
            end else if (5'h9 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_9;
            end else if (5'h8 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_8;
            end else if (5'h7 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_7;
            end else if (5'h6 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_6;
            end else if (5'h5 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_5;
            end else if (5'h4 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_4;
            end else if (5'h3 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_3;
            end else if (5'h2 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_2;
            end else if (5'h1 == _T_290[4:0]) begin
              rightNodeIsCharacter_0 <= isCharacter_1;
            end else begin
              rightNodeIsCharacter_0 <= isCharacter_0;
            end
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1 == validNodes[5:0]) begin
            if (5'h1f == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_31;
            end else if (5'h1e == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_30;
            end else if (5'h1d == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_29;
            end else if (5'h1c == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_28;
            end else if (5'h1b == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_27;
            end else if (5'h1a == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_26;
            end else if (5'h19 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_25;
            end else if (5'h18 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_24;
            end else if (5'h17 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_23;
            end else if (5'h16 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_22;
            end else if (5'h15 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_21;
            end else if (5'h14 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_20;
            end else if (5'h13 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_19;
            end else if (5'h12 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_18;
            end else if (5'h11 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_17;
            end else if (5'h10 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_16;
            end else if (5'hf == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_15;
            end else if (5'he == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_14;
            end else if (5'hd == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_13;
            end else if (5'hc == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_12;
            end else if (5'hb == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_11;
            end else if (5'ha == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_10;
            end else if (5'h9 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_9;
            end else if (5'h8 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_8;
            end else if (5'h7 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_7;
            end else if (5'h6 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_6;
            end else if (5'h5 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_5;
            end else if (5'h4 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_4;
            end else if (5'h3 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_3;
            end else if (5'h2 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_2;
            end else if (5'h1 == _T_290[4:0]) begin
              rightNodeIsCharacter_1 <= isCharacter_1;
            end else begin
              rightNodeIsCharacter_1 <= isCharacter_0;
            end
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2 == validNodes[5:0]) begin
            if (5'h1f == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_31;
            end else if (5'h1e == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_30;
            end else if (5'h1d == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_29;
            end else if (5'h1c == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_28;
            end else if (5'h1b == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_27;
            end else if (5'h1a == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_26;
            end else if (5'h19 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_25;
            end else if (5'h18 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_24;
            end else if (5'h17 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_23;
            end else if (5'h16 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_22;
            end else if (5'h15 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_21;
            end else if (5'h14 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_20;
            end else if (5'h13 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_19;
            end else if (5'h12 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_18;
            end else if (5'h11 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_17;
            end else if (5'h10 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_16;
            end else if (5'hf == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_15;
            end else if (5'he == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_14;
            end else if (5'hd == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_13;
            end else if (5'hc == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_12;
            end else if (5'hb == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_11;
            end else if (5'ha == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_10;
            end else if (5'h9 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_9;
            end else if (5'h8 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_8;
            end else if (5'h7 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_7;
            end else if (5'h6 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_6;
            end else if (5'h5 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_5;
            end else if (5'h4 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_4;
            end else if (5'h3 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_3;
            end else if (5'h2 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_2;
            end else if (5'h1 == _T_290[4:0]) begin
              rightNodeIsCharacter_2 <= isCharacter_1;
            end else begin
              rightNodeIsCharacter_2 <= isCharacter_0;
            end
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3 == validNodes[5:0]) begin
            if (5'h1f == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_31;
            end else if (5'h1e == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_30;
            end else if (5'h1d == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_29;
            end else if (5'h1c == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_28;
            end else if (5'h1b == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_27;
            end else if (5'h1a == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_26;
            end else if (5'h19 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_25;
            end else if (5'h18 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_24;
            end else if (5'h17 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_23;
            end else if (5'h16 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_22;
            end else if (5'h15 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_21;
            end else if (5'h14 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_20;
            end else if (5'h13 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_19;
            end else if (5'h12 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_18;
            end else if (5'h11 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_17;
            end else if (5'h10 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_16;
            end else if (5'hf == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_15;
            end else if (5'he == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_14;
            end else if (5'hd == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_13;
            end else if (5'hc == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_12;
            end else if (5'hb == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_11;
            end else if (5'ha == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_10;
            end else if (5'h9 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_9;
            end else if (5'h8 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_8;
            end else if (5'h7 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_7;
            end else if (5'h6 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_6;
            end else if (5'h5 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_5;
            end else if (5'h4 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_4;
            end else if (5'h3 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_3;
            end else if (5'h2 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_2;
            end else if (5'h1 == _T_290[4:0]) begin
              rightNodeIsCharacter_3 <= isCharacter_1;
            end else begin
              rightNodeIsCharacter_3 <= isCharacter_0;
            end
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h4 == validNodes[5:0]) begin
            rightNodeIsCharacter_4 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h5 == validNodes[5:0]) begin
            rightNodeIsCharacter_5 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h6 == validNodes[5:0]) begin
            rightNodeIsCharacter_6 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h7 == validNodes[5:0]) begin
            rightNodeIsCharacter_7 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h8 == validNodes[5:0]) begin
            rightNodeIsCharacter_8 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h9 == validNodes[5:0]) begin
            rightNodeIsCharacter_9 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'ha == validNodes[5:0]) begin
            rightNodeIsCharacter_10 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'hb == validNodes[5:0]) begin
            rightNodeIsCharacter_11 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'hc == validNodes[5:0]) begin
            rightNodeIsCharacter_12 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'hd == validNodes[5:0]) begin
            rightNodeIsCharacter_13 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'he == validNodes[5:0]) begin
            rightNodeIsCharacter_14 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'hf == validNodes[5:0]) begin
            rightNodeIsCharacter_15 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h10 == validNodes[5:0]) begin
            rightNodeIsCharacter_16 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h11 == validNodes[5:0]) begin
            rightNodeIsCharacter_17 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h12 == validNodes[5:0]) begin
            rightNodeIsCharacter_18 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h13 == validNodes[5:0]) begin
            rightNodeIsCharacter_19 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h14 == validNodes[5:0]) begin
            rightNodeIsCharacter_20 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h15 == validNodes[5:0]) begin
            rightNodeIsCharacter_21 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h16 == validNodes[5:0]) begin
            rightNodeIsCharacter_22 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h17 == validNodes[5:0]) begin
            rightNodeIsCharacter_23 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h18 == validNodes[5:0]) begin
            rightNodeIsCharacter_24 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h19 == validNodes[5:0]) begin
            rightNodeIsCharacter_25 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1a == validNodes[5:0]) begin
            rightNodeIsCharacter_26 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1b == validNodes[5:0]) begin
            rightNodeIsCharacter_27 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1c == validNodes[5:0]) begin
            rightNodeIsCharacter_28 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1d == validNodes[5:0]) begin
            rightNodeIsCharacter_29 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1e == validNodes[5:0]) begin
            rightNodeIsCharacter_30 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h1f == validNodes[5:0]) begin
            rightNodeIsCharacter_31 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h20 == validNodes[5:0]) begin
            rightNodeIsCharacter_32 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h21 == validNodes[5:0]) begin
            rightNodeIsCharacter_33 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h22 == validNodes[5:0]) begin
            rightNodeIsCharacter_34 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h23 == validNodes[5:0]) begin
            rightNodeIsCharacter_35 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h24 == validNodes[5:0]) begin
            rightNodeIsCharacter_36 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h25 == validNodes[5:0]) begin
            rightNodeIsCharacter_37 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h26 == validNodes[5:0]) begin
            rightNodeIsCharacter_38 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h27 == validNodes[5:0]) begin
            rightNodeIsCharacter_39 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h28 == validNodes[5:0]) begin
            rightNodeIsCharacter_40 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h29 == validNodes[5:0]) begin
            rightNodeIsCharacter_41 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2a == validNodes[5:0]) begin
            rightNodeIsCharacter_42 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2b == validNodes[5:0]) begin
            rightNodeIsCharacter_43 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2c == validNodes[5:0]) begin
            rightNodeIsCharacter_44 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2d == validNodes[5:0]) begin
            rightNodeIsCharacter_45 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2e == validNodes[5:0]) begin
            rightNodeIsCharacter_46 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h2f == validNodes[5:0]) begin
            rightNodeIsCharacter_47 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h30 == validNodes[5:0]) begin
            rightNodeIsCharacter_48 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h31 == validNodes[5:0]) begin
            rightNodeIsCharacter_49 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h32 == validNodes[5:0]) begin
            rightNodeIsCharacter_50 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h33 == validNodes[5:0]) begin
            rightNodeIsCharacter_51 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h34 == validNodes[5:0]) begin
            rightNodeIsCharacter_52 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h35 == validNodes[5:0]) begin
            rightNodeIsCharacter_53 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h36 == validNodes[5:0]) begin
            rightNodeIsCharacter_54 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h37 == validNodes[5:0]) begin
            rightNodeIsCharacter_55 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h38 == validNodes[5:0]) begin
            rightNodeIsCharacter_56 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h39 == validNodes[5:0]) begin
            rightNodeIsCharacter_57 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3a == validNodes[5:0]) begin
            rightNodeIsCharacter_58 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3b == validNodes[5:0]) begin
            rightNodeIsCharacter_59 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3c == validNodes[5:0]) begin
            rightNodeIsCharacter_60 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3d == validNodes[5:0]) begin
            rightNodeIsCharacter_61 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3e == validNodes[5:0]) begin
            rightNodeIsCharacter_62 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          if (6'h3f == validNodes[5:0]) begin
            rightNodeIsCharacter_63 <= _GEN_487;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          upperNodeIndex <= 6'h0;
        end
      end else if (_T_317) begin
        if (!(searchCompleted)) begin
          if (!(_T_404)) begin
            upperNodeIndex <= _T_402;
          end
        end
      end
    end
    if (!(_T_32)) begin
      if (_T_284) begin
        if (!(_T_285)) begin
          lowerNodeIndex <= _T_293;
        end
      end else if (_T_317) begin
        if (!(searchCompleted)) begin
          if (_T_404) begin
            lowerNodeIndex <= _T_402;
          end
        end
      end
    end
    if (_T_32) begin
      if (io_start) begin
        validNodes <= 7'h0;
      end
    end else if (_T_284) begin
      if (_T_285) begin
        if (_T_286) begin
          validNodes <= 7'h1;
        end
      end else begin
        validNodes <= _T_288;
      end
    end
    if (_T_32) begin
      if (io_start) begin
        validCharacters <= _T_157;
      end
    end else if (_T_284) begin
      if (_T_285) begin
        if (_T_286) begin
          validCharacters <= 6'h1;
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_32) begin
      if (io_start) begin
        state <= 2'h1;
      end
    end else if (_T_284) begin
      if (_T_285) begin
        state <= 2'h0;
      end else begin
        state <= 2'h2;
      end
    end else if (_T_317) begin
      if (searchCompleted) begin
        state <= 2'h1;
      end
    end
  end
endmodule
module treePathComparator(
  input  [31:0] io_position,
  input  [31:0] io_lastNode,
  input  [5:0]  io_length,
  output        io_equal
);
  wire [31:0] xorInputs = io_position ^ io_lastNode; // @[treePathComparator.scala 28:28]
  wire [31:0] _T_4 = {{16'd0}, xorInputs[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_6 = {xorInputs[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_8 = _T_6 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_9 = _T_4 | _T_8; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_0 = {{8'd0}, _T_9[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_14 = _GEN_0 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_16 = {_T_9[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_18 = _T_16 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_19 = _T_14 | _T_18; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1 = {{4'd0}, _T_19[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_24 = _GEN_1 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_26 = {_T_19[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_28 = _T_26 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_29 = _T_24 | _T_28; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_2 = {{2'd0}, _T_29[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_34 = _GEN_2 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_36 = {_T_29[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_38 = _T_36 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_39 = _T_34 | _T_38; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_3 = {{1'd0}, _T_39[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_44 = _GEN_3 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_46 = {_T_39[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_48 = _T_46 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire [31:0] _T_49 = _T_44 | _T_48; // @[Bitwise.scala 103:39]
  wire [32:0] reverseXor = {1'h1,_T_49}; // @[Cat.scala 29:58]
  wire [5:0] _T_84 = reverseXor[31] ? 6'h1f : 6'h20; // @[Mux.scala 47:69]
  wire [5:0] _T_85 = reverseXor[30] ? 6'h1e : _T_84; // @[Mux.scala 47:69]
  wire [5:0] _T_86 = reverseXor[29] ? 6'h1d : _T_85; // @[Mux.scala 47:69]
  wire [5:0] _T_87 = reverseXor[28] ? 6'h1c : _T_86; // @[Mux.scala 47:69]
  wire [5:0] _T_88 = reverseXor[27] ? 6'h1b : _T_87; // @[Mux.scala 47:69]
  wire [5:0] _T_89 = reverseXor[26] ? 6'h1a : _T_88; // @[Mux.scala 47:69]
  wire [5:0] _T_90 = reverseXor[25] ? 6'h19 : _T_89; // @[Mux.scala 47:69]
  wire [5:0] _T_91 = reverseXor[24] ? 6'h18 : _T_90; // @[Mux.scala 47:69]
  wire [5:0] _T_92 = reverseXor[23] ? 6'h17 : _T_91; // @[Mux.scala 47:69]
  wire [5:0] _T_93 = reverseXor[22] ? 6'h16 : _T_92; // @[Mux.scala 47:69]
  wire [5:0] _T_94 = reverseXor[21] ? 6'h15 : _T_93; // @[Mux.scala 47:69]
  wire [5:0] _T_95 = reverseXor[20] ? 6'h14 : _T_94; // @[Mux.scala 47:69]
  wire [5:0] _T_96 = reverseXor[19] ? 6'h13 : _T_95; // @[Mux.scala 47:69]
  wire [5:0] _T_97 = reverseXor[18] ? 6'h12 : _T_96; // @[Mux.scala 47:69]
  wire [5:0] _T_98 = reverseXor[17] ? 6'h11 : _T_97; // @[Mux.scala 47:69]
  wire [5:0] _T_99 = reverseXor[16] ? 6'h10 : _T_98; // @[Mux.scala 47:69]
  wire [5:0] _T_100 = reverseXor[15] ? 6'hf : _T_99; // @[Mux.scala 47:69]
  wire [5:0] _T_101 = reverseXor[14] ? 6'he : _T_100; // @[Mux.scala 47:69]
  wire [5:0] _T_102 = reverseXor[13] ? 6'hd : _T_101; // @[Mux.scala 47:69]
  wire [5:0] _T_103 = reverseXor[12] ? 6'hc : _T_102; // @[Mux.scala 47:69]
  wire [5:0] _T_104 = reverseXor[11] ? 6'hb : _T_103; // @[Mux.scala 47:69]
  wire [5:0] _T_105 = reverseXor[10] ? 6'ha : _T_104; // @[Mux.scala 47:69]
  wire [5:0] _T_106 = reverseXor[9] ? 6'h9 : _T_105; // @[Mux.scala 47:69]
  wire [5:0] _T_107 = reverseXor[8] ? 6'h8 : _T_106; // @[Mux.scala 47:69]
  wire [5:0] _T_108 = reverseXor[7] ? 6'h7 : _T_107; // @[Mux.scala 47:69]
  wire [5:0] _T_109 = reverseXor[6] ? 6'h6 : _T_108; // @[Mux.scala 47:69]
  wire [5:0] _T_110 = reverseXor[5] ? 6'h5 : _T_109; // @[Mux.scala 47:69]
  wire [5:0] _T_111 = reverseXor[4] ? 6'h4 : _T_110; // @[Mux.scala 47:69]
  wire [5:0] _T_112 = reverseXor[3] ? 6'h3 : _T_111; // @[Mux.scala 47:69]
  wire [5:0] _T_113 = reverseXor[2] ? 6'h2 : _T_112; // @[Mux.scala 47:69]
  wire [5:0] _T_114 = reverseXor[1] ? 6'h1 : _T_113; // @[Mux.scala 47:69]
  wire [5:0] _T_115 = reverseXor[0] ? 6'h0 : _T_114; // @[Mux.scala 47:69]
  assign io_equal = _T_115 >= io_length; // @[treePathComparator.scala 34:12]
endmodule
module treeDepthCounter(
  input        clock,
  input        reset,
  input        io_start,
  input  [8:0] io_inputs_leftNode_0,
  input  [8:0] io_inputs_leftNode_1,
  input  [8:0] io_inputs_leftNode_2,
  input  [8:0] io_inputs_leftNode_3,
  input  [8:0] io_inputs_leftNode_4,
  input  [8:0] io_inputs_leftNode_5,
  input  [8:0] io_inputs_leftNode_6,
  input  [8:0] io_inputs_leftNode_7,
  input  [8:0] io_inputs_leftNode_8,
  input  [8:0] io_inputs_leftNode_9,
  input  [8:0] io_inputs_leftNode_10,
  input  [8:0] io_inputs_leftNode_11,
  input  [8:0] io_inputs_leftNode_12,
  input  [8:0] io_inputs_leftNode_13,
  input  [8:0] io_inputs_leftNode_14,
  input  [8:0] io_inputs_leftNode_15,
  input  [8:0] io_inputs_leftNode_16,
  input  [8:0] io_inputs_leftNode_17,
  input  [8:0] io_inputs_leftNode_18,
  input  [8:0] io_inputs_leftNode_19,
  input  [8:0] io_inputs_leftNode_20,
  input  [8:0] io_inputs_leftNode_21,
  input  [8:0] io_inputs_leftNode_22,
  input  [8:0] io_inputs_leftNode_23,
  input  [8:0] io_inputs_leftNode_24,
  input  [8:0] io_inputs_leftNode_25,
  input  [8:0] io_inputs_leftNode_26,
  input  [8:0] io_inputs_leftNode_27,
  input  [8:0] io_inputs_leftNode_28,
  input  [8:0] io_inputs_leftNode_29,
  input  [8:0] io_inputs_leftNode_30,
  input  [8:0] io_inputs_leftNode_31,
  input  [8:0] io_inputs_leftNode_32,
  input  [8:0] io_inputs_leftNode_33,
  input  [8:0] io_inputs_leftNode_34,
  input  [8:0] io_inputs_leftNode_35,
  input  [8:0] io_inputs_leftNode_36,
  input  [8:0] io_inputs_leftNode_37,
  input  [8:0] io_inputs_leftNode_38,
  input  [8:0] io_inputs_leftNode_39,
  input  [8:0] io_inputs_leftNode_40,
  input  [8:0] io_inputs_leftNode_41,
  input  [8:0] io_inputs_leftNode_42,
  input  [8:0] io_inputs_leftNode_43,
  input  [8:0] io_inputs_leftNode_44,
  input  [8:0] io_inputs_leftNode_45,
  input  [8:0] io_inputs_leftNode_46,
  input  [8:0] io_inputs_leftNode_47,
  input  [8:0] io_inputs_leftNode_48,
  input  [8:0] io_inputs_leftNode_49,
  input  [8:0] io_inputs_leftNode_50,
  input  [8:0] io_inputs_leftNode_51,
  input  [8:0] io_inputs_leftNode_52,
  input  [8:0] io_inputs_leftNode_53,
  input  [8:0] io_inputs_leftNode_54,
  input  [8:0] io_inputs_leftNode_55,
  input  [8:0] io_inputs_leftNode_56,
  input  [8:0] io_inputs_leftNode_57,
  input  [8:0] io_inputs_leftNode_58,
  input  [8:0] io_inputs_leftNode_59,
  input  [8:0] io_inputs_leftNode_60,
  input  [8:0] io_inputs_leftNode_61,
  input  [8:0] io_inputs_leftNode_62,
  input  [8:0] io_inputs_leftNode_63,
  input  [8:0] io_inputs_rightNode_0,
  input  [8:0] io_inputs_rightNode_1,
  input  [8:0] io_inputs_rightNode_2,
  input  [8:0] io_inputs_rightNode_3,
  input  [8:0] io_inputs_rightNode_4,
  input  [8:0] io_inputs_rightNode_5,
  input  [8:0] io_inputs_rightNode_6,
  input  [8:0] io_inputs_rightNode_7,
  input  [8:0] io_inputs_rightNode_8,
  input  [8:0] io_inputs_rightNode_9,
  input  [8:0] io_inputs_rightNode_10,
  input  [8:0] io_inputs_rightNode_11,
  input  [8:0] io_inputs_rightNode_12,
  input  [8:0] io_inputs_rightNode_13,
  input  [8:0] io_inputs_rightNode_14,
  input  [8:0] io_inputs_rightNode_15,
  input  [8:0] io_inputs_rightNode_16,
  input  [8:0] io_inputs_rightNode_17,
  input  [8:0] io_inputs_rightNode_18,
  input  [8:0] io_inputs_rightNode_19,
  input  [8:0] io_inputs_rightNode_20,
  input  [8:0] io_inputs_rightNode_21,
  input  [8:0] io_inputs_rightNode_22,
  input  [8:0] io_inputs_rightNode_23,
  input  [8:0] io_inputs_rightNode_24,
  input  [8:0] io_inputs_rightNode_25,
  input  [8:0] io_inputs_rightNode_26,
  input  [8:0] io_inputs_rightNode_27,
  input  [8:0] io_inputs_rightNode_28,
  input  [8:0] io_inputs_rightNode_29,
  input  [8:0] io_inputs_rightNode_30,
  input  [8:0] io_inputs_rightNode_31,
  input  [8:0] io_inputs_rightNode_32,
  input  [8:0] io_inputs_rightNode_33,
  input  [8:0] io_inputs_rightNode_34,
  input  [8:0] io_inputs_rightNode_35,
  input  [8:0] io_inputs_rightNode_36,
  input  [8:0] io_inputs_rightNode_37,
  input  [8:0] io_inputs_rightNode_38,
  input  [8:0] io_inputs_rightNode_39,
  input  [8:0] io_inputs_rightNode_40,
  input  [8:0] io_inputs_rightNode_41,
  input  [8:0] io_inputs_rightNode_42,
  input  [8:0] io_inputs_rightNode_43,
  input  [8:0] io_inputs_rightNode_44,
  input  [8:0] io_inputs_rightNode_45,
  input  [8:0] io_inputs_rightNode_46,
  input  [8:0] io_inputs_rightNode_47,
  input  [8:0] io_inputs_rightNode_48,
  input  [8:0] io_inputs_rightNode_49,
  input  [8:0] io_inputs_rightNode_50,
  input  [8:0] io_inputs_rightNode_51,
  input  [8:0] io_inputs_rightNode_52,
  input  [8:0] io_inputs_rightNode_53,
  input  [8:0] io_inputs_rightNode_54,
  input  [8:0] io_inputs_rightNode_55,
  input  [8:0] io_inputs_rightNode_56,
  input  [8:0] io_inputs_rightNode_57,
  input  [8:0] io_inputs_rightNode_58,
  input  [8:0] io_inputs_rightNode_59,
  input  [8:0] io_inputs_rightNode_60,
  input  [8:0] io_inputs_rightNode_61,
  input  [8:0] io_inputs_rightNode_62,
  input  [8:0] io_inputs_rightNode_63,
  input        io_inputs_leftNodeIsCharacter_0,
  input        io_inputs_leftNodeIsCharacter_1,
  input        io_inputs_leftNodeIsCharacter_2,
  input        io_inputs_leftNodeIsCharacter_3,
  input        io_inputs_leftNodeIsCharacter_4,
  input        io_inputs_leftNodeIsCharacter_5,
  input        io_inputs_leftNodeIsCharacter_6,
  input        io_inputs_leftNodeIsCharacter_7,
  input        io_inputs_leftNodeIsCharacter_8,
  input        io_inputs_leftNodeIsCharacter_9,
  input        io_inputs_leftNodeIsCharacter_10,
  input        io_inputs_leftNodeIsCharacter_11,
  input        io_inputs_leftNodeIsCharacter_12,
  input        io_inputs_leftNodeIsCharacter_13,
  input        io_inputs_leftNodeIsCharacter_14,
  input        io_inputs_leftNodeIsCharacter_15,
  input        io_inputs_leftNodeIsCharacter_16,
  input        io_inputs_leftNodeIsCharacter_17,
  input        io_inputs_leftNodeIsCharacter_18,
  input        io_inputs_leftNodeIsCharacter_19,
  input        io_inputs_leftNodeIsCharacter_20,
  input        io_inputs_leftNodeIsCharacter_21,
  input        io_inputs_leftNodeIsCharacter_22,
  input        io_inputs_leftNodeIsCharacter_23,
  input        io_inputs_leftNodeIsCharacter_24,
  input        io_inputs_leftNodeIsCharacter_25,
  input        io_inputs_leftNodeIsCharacter_26,
  input        io_inputs_leftNodeIsCharacter_27,
  input        io_inputs_leftNodeIsCharacter_28,
  input        io_inputs_leftNodeIsCharacter_29,
  input        io_inputs_leftNodeIsCharacter_30,
  input        io_inputs_leftNodeIsCharacter_31,
  input        io_inputs_leftNodeIsCharacter_32,
  input        io_inputs_leftNodeIsCharacter_33,
  input        io_inputs_leftNodeIsCharacter_34,
  input        io_inputs_leftNodeIsCharacter_35,
  input        io_inputs_leftNodeIsCharacter_36,
  input        io_inputs_leftNodeIsCharacter_37,
  input        io_inputs_leftNodeIsCharacter_38,
  input        io_inputs_leftNodeIsCharacter_39,
  input        io_inputs_leftNodeIsCharacter_40,
  input        io_inputs_leftNodeIsCharacter_41,
  input        io_inputs_leftNodeIsCharacter_42,
  input        io_inputs_leftNodeIsCharacter_43,
  input        io_inputs_leftNodeIsCharacter_44,
  input        io_inputs_leftNodeIsCharacter_45,
  input        io_inputs_leftNodeIsCharacter_46,
  input        io_inputs_leftNodeIsCharacter_47,
  input        io_inputs_leftNodeIsCharacter_48,
  input        io_inputs_leftNodeIsCharacter_49,
  input        io_inputs_leftNodeIsCharacter_50,
  input        io_inputs_leftNodeIsCharacter_51,
  input        io_inputs_leftNodeIsCharacter_52,
  input        io_inputs_leftNodeIsCharacter_53,
  input        io_inputs_leftNodeIsCharacter_54,
  input        io_inputs_leftNodeIsCharacter_55,
  input        io_inputs_leftNodeIsCharacter_56,
  input        io_inputs_leftNodeIsCharacter_57,
  input        io_inputs_leftNodeIsCharacter_58,
  input        io_inputs_leftNodeIsCharacter_59,
  input        io_inputs_leftNodeIsCharacter_60,
  input        io_inputs_leftNodeIsCharacter_61,
  input        io_inputs_leftNodeIsCharacter_62,
  input        io_inputs_leftNodeIsCharacter_63,
  input        io_inputs_rightNodeIsCharacter_0,
  input        io_inputs_rightNodeIsCharacter_1,
  input        io_inputs_rightNodeIsCharacter_2,
  input        io_inputs_rightNodeIsCharacter_3,
  input        io_inputs_rightNodeIsCharacter_4,
  input        io_inputs_rightNodeIsCharacter_5,
  input        io_inputs_rightNodeIsCharacter_6,
  input        io_inputs_rightNodeIsCharacter_7,
  input        io_inputs_rightNodeIsCharacter_8,
  input        io_inputs_rightNodeIsCharacter_9,
  input        io_inputs_rightNodeIsCharacter_10,
  input        io_inputs_rightNodeIsCharacter_11,
  input        io_inputs_rightNodeIsCharacter_12,
  input        io_inputs_rightNodeIsCharacter_13,
  input        io_inputs_rightNodeIsCharacter_14,
  input        io_inputs_rightNodeIsCharacter_15,
  input        io_inputs_rightNodeIsCharacter_16,
  input        io_inputs_rightNodeIsCharacter_17,
  input        io_inputs_rightNodeIsCharacter_18,
  input        io_inputs_rightNodeIsCharacter_19,
  input        io_inputs_rightNodeIsCharacter_20,
  input        io_inputs_rightNodeIsCharacter_21,
  input        io_inputs_rightNodeIsCharacter_22,
  input        io_inputs_rightNodeIsCharacter_23,
  input        io_inputs_rightNodeIsCharacter_24,
  input        io_inputs_rightNodeIsCharacter_25,
  input        io_inputs_rightNodeIsCharacter_26,
  input        io_inputs_rightNodeIsCharacter_27,
  input        io_inputs_rightNodeIsCharacter_28,
  input        io_inputs_rightNodeIsCharacter_29,
  input        io_inputs_rightNodeIsCharacter_30,
  input        io_inputs_rightNodeIsCharacter_31,
  input        io_inputs_rightNodeIsCharacter_32,
  input        io_inputs_rightNodeIsCharacter_33,
  input        io_inputs_rightNodeIsCharacter_34,
  input        io_inputs_rightNodeIsCharacter_35,
  input        io_inputs_rightNodeIsCharacter_36,
  input        io_inputs_rightNodeIsCharacter_37,
  input        io_inputs_rightNodeIsCharacter_38,
  input        io_inputs_rightNodeIsCharacter_39,
  input        io_inputs_rightNodeIsCharacter_40,
  input        io_inputs_rightNodeIsCharacter_41,
  input        io_inputs_rightNodeIsCharacter_42,
  input        io_inputs_rightNodeIsCharacter_43,
  input        io_inputs_rightNodeIsCharacter_44,
  input        io_inputs_rightNodeIsCharacter_45,
  input        io_inputs_rightNodeIsCharacter_46,
  input        io_inputs_rightNodeIsCharacter_47,
  input        io_inputs_rightNodeIsCharacter_48,
  input        io_inputs_rightNodeIsCharacter_49,
  input        io_inputs_rightNodeIsCharacter_50,
  input        io_inputs_rightNodeIsCharacter_51,
  input        io_inputs_rightNodeIsCharacter_52,
  input        io_inputs_rightNodeIsCharacter_53,
  input        io_inputs_rightNodeIsCharacter_54,
  input        io_inputs_rightNodeIsCharacter_55,
  input        io_inputs_rightNodeIsCharacter_56,
  input        io_inputs_rightNodeIsCharacter_57,
  input        io_inputs_rightNodeIsCharacter_58,
  input        io_inputs_rightNodeIsCharacter_59,
  input        io_inputs_rightNodeIsCharacter_60,
  input        io_inputs_rightNodeIsCharacter_61,
  input        io_inputs_rightNodeIsCharacter_62,
  input        io_inputs_rightNodeIsCharacter_63,
  input  [6:0] io_inputs_validNodes,
  input  [5:0] io_inputs_validCharacters,
  output [8:0] io_outputs_characters_0,
  output [8:0] io_outputs_characters_1,
  output [8:0] io_outputs_characters_2,
  output [8:0] io_outputs_characters_3,
  output [8:0] io_outputs_characters_4,
  output [8:0] io_outputs_characters_5,
  output [8:0] io_outputs_characters_6,
  output [8:0] io_outputs_characters_7,
  output [8:0] io_outputs_characters_8,
  output [8:0] io_outputs_characters_9,
  output [8:0] io_outputs_characters_10,
  output [8:0] io_outputs_characters_11,
  output [8:0] io_outputs_characters_12,
  output [8:0] io_outputs_characters_13,
  output [8:0] io_outputs_characters_14,
  output [8:0] io_outputs_characters_15,
  output [8:0] io_outputs_characters_16,
  output [8:0] io_outputs_characters_17,
  output [8:0] io_outputs_characters_18,
  output [8:0] io_outputs_characters_19,
  output [8:0] io_outputs_characters_20,
  output [8:0] io_outputs_characters_21,
  output [8:0] io_outputs_characters_22,
  output [8:0] io_outputs_characters_23,
  output [8:0] io_outputs_characters_24,
  output [8:0] io_outputs_characters_25,
  output [8:0] io_outputs_characters_26,
  output [8:0] io_outputs_characters_27,
  output [8:0] io_outputs_characters_28,
  output [8:0] io_outputs_characters_29,
  output [8:0] io_outputs_characters_30,
  output [8:0] io_outputs_characters_31,
  output [5:0] io_outputs_depths_0,
  output [5:0] io_outputs_depths_1,
  output [5:0] io_outputs_depths_2,
  output [5:0] io_outputs_depths_3,
  output [5:0] io_outputs_depths_4,
  output [5:0] io_outputs_depths_5,
  output [5:0] io_outputs_depths_6,
  output [5:0] io_outputs_depths_7,
  output [5:0] io_outputs_depths_8,
  output [5:0] io_outputs_depths_9,
  output [5:0] io_outputs_depths_10,
  output [5:0] io_outputs_depths_11,
  output [5:0] io_outputs_depths_12,
  output [5:0] io_outputs_depths_13,
  output [5:0] io_outputs_depths_14,
  output [5:0] io_outputs_depths_15,
  output [5:0] io_outputs_depths_16,
  output [5:0] io_outputs_depths_17,
  output [5:0] io_outputs_depths_18,
  output [5:0] io_outputs_depths_19,
  output [5:0] io_outputs_depths_20,
  output [5:0] io_outputs_depths_21,
  output [5:0] io_outputs_depths_22,
  output [5:0] io_outputs_depths_23,
  output [5:0] io_outputs_depths_24,
  output [5:0] io_outputs_depths_25,
  output [5:0] io_outputs_depths_26,
  output [5:0] io_outputs_depths_27,
  output [5:0] io_outputs_depths_28,
  output [5:0] io_outputs_depths_29,
  output [5:0] io_outputs_depths_30,
  output [5:0] io_outputs_depths_31,
  output [5:0] io_outputs_validCharacters,
  output       io_finished
);
  wire [31:0] tpc_io_position; // @[treeDepthCounter.scala 45:19]
  wire [31:0] tpc_io_lastNode; // @[treeDepthCounter.scala 45:19]
  wire [5:0] tpc_io_length; // @[treeDepthCounter.scala 45:19]
  wire  tpc_io_equal; // @[treeDepthCounter.scala 45:19]
  reg [8:0] leftNode_0; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_0;
  reg [8:0] leftNode_1; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_1;
  reg [8:0] leftNode_2; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_2;
  reg [8:0] leftNode_3; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_3;
  reg [8:0] leftNode_4; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_4;
  reg [8:0] leftNode_5; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_5;
  reg [8:0] leftNode_6; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_6;
  reg [8:0] leftNode_7; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_7;
  reg [8:0] leftNode_8; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_8;
  reg [8:0] leftNode_9; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_9;
  reg [8:0] leftNode_10; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_10;
  reg [8:0] leftNode_11; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_11;
  reg [8:0] leftNode_12; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_12;
  reg [8:0] leftNode_13; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_13;
  reg [8:0] leftNode_14; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_14;
  reg [8:0] leftNode_15; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_15;
  reg [8:0] leftNode_16; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_16;
  reg [8:0] leftNode_17; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_17;
  reg [8:0] leftNode_18; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_18;
  reg [8:0] leftNode_19; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_19;
  reg [8:0] leftNode_20; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_20;
  reg [8:0] leftNode_21; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_21;
  reg [8:0] leftNode_22; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_22;
  reg [8:0] leftNode_23; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_23;
  reg [8:0] leftNode_24; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_24;
  reg [8:0] leftNode_25; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_25;
  reg [8:0] leftNode_26; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_26;
  reg [8:0] leftNode_27; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_27;
  reg [8:0] leftNode_28; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_28;
  reg [8:0] leftNode_29; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_29;
  reg [8:0] leftNode_30; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_30;
  reg [8:0] leftNode_31; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_31;
  reg [8:0] leftNode_32; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_32;
  reg [8:0] leftNode_33; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_33;
  reg [8:0] leftNode_34; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_34;
  reg [8:0] leftNode_35; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_35;
  reg [8:0] leftNode_36; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_36;
  reg [8:0] leftNode_37; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_37;
  reg [8:0] leftNode_38; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_38;
  reg [8:0] leftNode_39; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_39;
  reg [8:0] leftNode_40; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_40;
  reg [8:0] leftNode_41; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_41;
  reg [8:0] leftNode_42; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_42;
  reg [8:0] leftNode_43; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_43;
  reg [8:0] leftNode_44; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_44;
  reg [8:0] leftNode_45; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_45;
  reg [8:0] leftNode_46; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_46;
  reg [8:0] leftNode_47; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_47;
  reg [8:0] leftNode_48; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_48;
  reg [8:0] leftNode_49; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_49;
  reg [8:0] leftNode_50; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_50;
  reg [8:0] leftNode_51; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_51;
  reg [8:0] leftNode_52; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_52;
  reg [8:0] leftNode_53; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_53;
  reg [8:0] leftNode_54; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_54;
  reg [8:0] leftNode_55; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_55;
  reg [8:0] leftNode_56; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_56;
  reg [8:0] leftNode_57; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_57;
  reg [8:0] leftNode_58; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_58;
  reg [8:0] leftNode_59; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_59;
  reg [8:0] leftNode_60; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_60;
  reg [8:0] leftNode_61; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_61;
  reg [8:0] leftNode_62; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_62;
  reg [8:0] leftNode_63; // @[treeDepthCounter.scala 18:21]
  reg [31:0] _RAND_63;
  reg [8:0] rightNode_0; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_64;
  reg [8:0] rightNode_1; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_65;
  reg [8:0] rightNode_2; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_66;
  reg [8:0] rightNode_3; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_67;
  reg [8:0] rightNode_4; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_68;
  reg [8:0] rightNode_5; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_69;
  reg [8:0] rightNode_6; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_70;
  reg [8:0] rightNode_7; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_71;
  reg [8:0] rightNode_8; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_72;
  reg [8:0] rightNode_9; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_73;
  reg [8:0] rightNode_10; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_74;
  reg [8:0] rightNode_11; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_75;
  reg [8:0] rightNode_12; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_76;
  reg [8:0] rightNode_13; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_77;
  reg [8:0] rightNode_14; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_78;
  reg [8:0] rightNode_15; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_79;
  reg [8:0] rightNode_16; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_80;
  reg [8:0] rightNode_17; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_81;
  reg [8:0] rightNode_18; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_82;
  reg [8:0] rightNode_19; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_83;
  reg [8:0] rightNode_20; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_84;
  reg [8:0] rightNode_21; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_85;
  reg [8:0] rightNode_22; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_86;
  reg [8:0] rightNode_23; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_87;
  reg [8:0] rightNode_24; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_88;
  reg [8:0] rightNode_25; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_89;
  reg [8:0] rightNode_26; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_90;
  reg [8:0] rightNode_27; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_91;
  reg [8:0] rightNode_28; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_92;
  reg [8:0] rightNode_29; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_93;
  reg [8:0] rightNode_30; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_94;
  reg [8:0] rightNode_31; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_95;
  reg [8:0] rightNode_32; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_96;
  reg [8:0] rightNode_33; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_97;
  reg [8:0] rightNode_34; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_98;
  reg [8:0] rightNode_35; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_99;
  reg [8:0] rightNode_36; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_100;
  reg [8:0] rightNode_37; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_101;
  reg [8:0] rightNode_38; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_102;
  reg [8:0] rightNode_39; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_103;
  reg [8:0] rightNode_40; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_104;
  reg [8:0] rightNode_41; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_105;
  reg [8:0] rightNode_42; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_106;
  reg [8:0] rightNode_43; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_107;
  reg [8:0] rightNode_44; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_108;
  reg [8:0] rightNode_45; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_109;
  reg [8:0] rightNode_46; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_110;
  reg [8:0] rightNode_47; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_111;
  reg [8:0] rightNode_48; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_112;
  reg [8:0] rightNode_49; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_113;
  reg [8:0] rightNode_50; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_114;
  reg [8:0] rightNode_51; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_115;
  reg [8:0] rightNode_52; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_116;
  reg [8:0] rightNode_53; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_117;
  reg [8:0] rightNode_54; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_118;
  reg [8:0] rightNode_55; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_119;
  reg [8:0] rightNode_56; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_120;
  reg [8:0] rightNode_57; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_121;
  reg [8:0] rightNode_58; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_122;
  reg [8:0] rightNode_59; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_123;
  reg [8:0] rightNode_60; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_124;
  reg [8:0] rightNode_61; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_125;
  reg [8:0] rightNode_62; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_126;
  reg [8:0] rightNode_63; // @[treeDepthCounter.scala 21:22]
  reg [31:0] _RAND_127;
  reg  leftNodeIsCharacter_0; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_128;
  reg  leftNodeIsCharacter_1; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_129;
  reg  leftNodeIsCharacter_2; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_130;
  reg  leftNodeIsCharacter_3; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_131;
  reg  leftNodeIsCharacter_4; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_132;
  reg  leftNodeIsCharacter_5; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_133;
  reg  leftNodeIsCharacter_6; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_134;
  reg  leftNodeIsCharacter_7; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_135;
  reg  leftNodeIsCharacter_8; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_136;
  reg  leftNodeIsCharacter_9; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_137;
  reg  leftNodeIsCharacter_10; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_138;
  reg  leftNodeIsCharacter_11; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_139;
  reg  leftNodeIsCharacter_12; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_140;
  reg  leftNodeIsCharacter_13; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_141;
  reg  leftNodeIsCharacter_14; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_142;
  reg  leftNodeIsCharacter_15; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_143;
  reg  leftNodeIsCharacter_16; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_144;
  reg  leftNodeIsCharacter_17; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_145;
  reg  leftNodeIsCharacter_18; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_146;
  reg  leftNodeIsCharacter_19; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_147;
  reg  leftNodeIsCharacter_20; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_148;
  reg  leftNodeIsCharacter_21; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_149;
  reg  leftNodeIsCharacter_22; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_150;
  reg  leftNodeIsCharacter_23; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_151;
  reg  leftNodeIsCharacter_24; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_152;
  reg  leftNodeIsCharacter_25; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_153;
  reg  leftNodeIsCharacter_26; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_154;
  reg  leftNodeIsCharacter_27; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_155;
  reg  leftNodeIsCharacter_28; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_156;
  reg  leftNodeIsCharacter_29; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_157;
  reg  leftNodeIsCharacter_30; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_158;
  reg  leftNodeIsCharacter_31; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_159;
  reg  leftNodeIsCharacter_32; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_160;
  reg  leftNodeIsCharacter_33; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_161;
  reg  leftNodeIsCharacter_34; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_162;
  reg  leftNodeIsCharacter_35; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_163;
  reg  leftNodeIsCharacter_36; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_164;
  reg  leftNodeIsCharacter_37; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_165;
  reg  leftNodeIsCharacter_38; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_166;
  reg  leftNodeIsCharacter_39; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_167;
  reg  leftNodeIsCharacter_40; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_168;
  reg  leftNodeIsCharacter_41; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_169;
  reg  leftNodeIsCharacter_42; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_170;
  reg  leftNodeIsCharacter_43; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_171;
  reg  leftNodeIsCharacter_44; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_172;
  reg  leftNodeIsCharacter_45; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_173;
  reg  leftNodeIsCharacter_46; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_174;
  reg  leftNodeIsCharacter_47; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_175;
  reg  leftNodeIsCharacter_48; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_176;
  reg  leftNodeIsCharacter_49; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_177;
  reg  leftNodeIsCharacter_50; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_178;
  reg  leftNodeIsCharacter_51; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_179;
  reg  leftNodeIsCharacter_52; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_180;
  reg  leftNodeIsCharacter_53; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_181;
  reg  leftNodeIsCharacter_54; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_182;
  reg  leftNodeIsCharacter_55; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_183;
  reg  leftNodeIsCharacter_56; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_184;
  reg  leftNodeIsCharacter_57; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_185;
  reg  leftNodeIsCharacter_58; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_186;
  reg  leftNodeIsCharacter_59; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_187;
  reg  leftNodeIsCharacter_60; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_188;
  reg  leftNodeIsCharacter_61; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_189;
  reg  leftNodeIsCharacter_62; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_190;
  reg  leftNodeIsCharacter_63; // @[treeDepthCounter.scala 24:32]
  reg [31:0] _RAND_191;
  reg  rightNodeIsCharacter_0; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_192;
  reg  rightNodeIsCharacter_1; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_193;
  reg  rightNodeIsCharacter_2; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_194;
  reg  rightNodeIsCharacter_3; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_195;
  reg  rightNodeIsCharacter_4; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_196;
  reg  rightNodeIsCharacter_5; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_197;
  reg  rightNodeIsCharacter_6; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_198;
  reg  rightNodeIsCharacter_7; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_199;
  reg  rightNodeIsCharacter_8; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_200;
  reg  rightNodeIsCharacter_9; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_201;
  reg  rightNodeIsCharacter_10; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_202;
  reg  rightNodeIsCharacter_11; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_203;
  reg  rightNodeIsCharacter_12; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_204;
  reg  rightNodeIsCharacter_13; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_205;
  reg  rightNodeIsCharacter_14; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_206;
  reg  rightNodeIsCharacter_15; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_207;
  reg  rightNodeIsCharacter_16; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_208;
  reg  rightNodeIsCharacter_17; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_209;
  reg  rightNodeIsCharacter_18; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_210;
  reg  rightNodeIsCharacter_19; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_211;
  reg  rightNodeIsCharacter_20; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_212;
  reg  rightNodeIsCharacter_21; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_213;
  reg  rightNodeIsCharacter_22; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_214;
  reg  rightNodeIsCharacter_23; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_215;
  reg  rightNodeIsCharacter_24; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_216;
  reg  rightNodeIsCharacter_25; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_217;
  reg  rightNodeIsCharacter_26; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_218;
  reg  rightNodeIsCharacter_27; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_219;
  reg  rightNodeIsCharacter_28; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_220;
  reg  rightNodeIsCharacter_29; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_221;
  reg  rightNodeIsCharacter_30; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_222;
  reg  rightNodeIsCharacter_31; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_223;
  reg  rightNodeIsCharacter_32; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_224;
  reg  rightNodeIsCharacter_33; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_225;
  reg  rightNodeIsCharacter_34; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_226;
  reg  rightNodeIsCharacter_35; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_227;
  reg  rightNodeIsCharacter_36; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_228;
  reg  rightNodeIsCharacter_37; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_229;
  reg  rightNodeIsCharacter_38; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_230;
  reg  rightNodeIsCharacter_39; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_231;
  reg  rightNodeIsCharacter_40; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_232;
  reg  rightNodeIsCharacter_41; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_233;
  reg  rightNodeIsCharacter_42; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_234;
  reg  rightNodeIsCharacter_43; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_235;
  reg  rightNodeIsCharacter_44; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_236;
  reg  rightNodeIsCharacter_45; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_237;
  reg  rightNodeIsCharacter_46; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_238;
  reg  rightNodeIsCharacter_47; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_239;
  reg  rightNodeIsCharacter_48; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_240;
  reg  rightNodeIsCharacter_49; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_241;
  reg  rightNodeIsCharacter_50; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_242;
  reg  rightNodeIsCharacter_51; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_243;
  reg  rightNodeIsCharacter_52; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_244;
  reg  rightNodeIsCharacter_53; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_245;
  reg  rightNodeIsCharacter_54; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_246;
  reg  rightNodeIsCharacter_55; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_247;
  reg  rightNodeIsCharacter_56; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_248;
  reg  rightNodeIsCharacter_57; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_249;
  reg  rightNodeIsCharacter_58; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_250;
  reg  rightNodeIsCharacter_59; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_251;
  reg  rightNodeIsCharacter_60; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_252;
  reg  rightNodeIsCharacter_61; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_253;
  reg  rightNodeIsCharacter_62; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_254;
  reg  rightNodeIsCharacter_63; // @[treeDepthCounter.scala 25:33]
  reg [31:0] _RAND_255;
  reg [5:0] validCharacters; // @[treeDepthCounter.scala 26:28]
  reg [31:0] _RAND_256;
  reg [5:0] charactersVisited; // @[treeDepthCounter.scala 28:30]
  reg [31:0] _RAND_257;
  reg [8:0] parentNodes_0; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_258;
  reg [8:0] parentNodes_1; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_259;
  reg [8:0] parentNodes_2; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_260;
  reg [8:0] parentNodes_3; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_261;
  reg [8:0] parentNodes_4; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_262;
  reg [8:0] parentNodes_5; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_263;
  reg [8:0] parentNodes_6; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_264;
  reg [8:0] parentNodes_7; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_265;
  reg [8:0] parentNodes_8; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_266;
  reg [8:0] parentNodes_9; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_267;
  reg [8:0] parentNodes_10; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_268;
  reg [8:0] parentNodes_11; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_269;
  reg [8:0] parentNodes_12; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_270;
  reg [8:0] parentNodes_13; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_271;
  reg [8:0] parentNodes_14; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_272;
  reg [8:0] parentNodes_15; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_273;
  reg [8:0] parentNodes_16; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_274;
  reg [8:0] parentNodes_17; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_275;
  reg [8:0] parentNodes_18; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_276;
  reg [8:0] parentNodes_19; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_277;
  reg [8:0] parentNodes_20; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_278;
  reg [8:0] parentNodes_21; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_279;
  reg [8:0] parentNodes_22; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_280;
  reg [8:0] parentNodes_23; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_281;
  reg [8:0] parentNodes_24; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_282;
  reg [8:0] parentNodes_25; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_283;
  reg [8:0] parentNodes_26; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_284;
  reg [8:0] parentNodes_27; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_285;
  reg [8:0] parentNodes_28; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_286;
  reg [8:0] parentNodes_29; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_287;
  reg [8:0] parentNodes_30; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_288;
  reg [8:0] parentNodes_31; // @[treeDepthCounter.scala 30:24]
  reg [31:0] _RAND_289;
  reg [31:0] position; // @[treeDepthCounter.scala 39:21]
  reg [31:0] _RAND_290;
  reg [31:0] lastNode; // @[treeDepthCounter.scala 40:21]
  reg [31:0] _RAND_291;
  reg [5:0] positionDepth; // @[treeDepthCounter.scala 41:26]
  reg [31:0] _RAND_292;
  reg [5:0] lastNodeDepth; // @[treeDepthCounter.scala 42:26]
  reg [31:0] _RAND_293;
  reg [8:0] characters_0; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_294;
  reg [8:0] characters_1; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_295;
  reg [8:0] characters_2; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_296;
  reg [8:0] characters_3; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_297;
  reg [8:0] characters_4; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_298;
  reg [8:0] characters_5; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_299;
  reg [8:0] characters_6; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_300;
  reg [8:0] characters_7; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_301;
  reg [8:0] characters_8; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_302;
  reg [8:0] characters_9; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_303;
  reg [8:0] characters_10; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_304;
  reg [8:0] characters_11; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_305;
  reg [8:0] characters_12; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_306;
  reg [8:0] characters_13; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_307;
  reg [8:0] characters_14; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_308;
  reg [8:0] characters_15; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_309;
  reg [8:0] characters_16; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_310;
  reg [8:0] characters_17; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_311;
  reg [8:0] characters_18; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_312;
  reg [8:0] characters_19; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_313;
  reg [8:0] characters_20; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_314;
  reg [8:0] characters_21; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_315;
  reg [8:0] characters_22; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_316;
  reg [8:0] characters_23; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_317;
  reg [8:0] characters_24; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_318;
  reg [8:0] characters_25; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_319;
  reg [8:0] characters_26; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_320;
  reg [8:0] characters_27; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_321;
  reg [8:0] characters_28; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_322;
  reg [8:0] characters_29; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_323;
  reg [8:0] characters_30; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_324;
  reg [8:0] characters_31; // @[treeDepthCounter.scala 50:23]
  reg [31:0] _RAND_325;
  reg [5:0] depths_0; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_326;
  reg [5:0] depths_1; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_327;
  reg [5:0] depths_2; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_328;
  reg [5:0] depths_3; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_329;
  reg [5:0] depths_4; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_330;
  reg [5:0] depths_5; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_331;
  reg [5:0] depths_6; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_332;
  reg [5:0] depths_7; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_333;
  reg [5:0] depths_8; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_334;
  reg [5:0] depths_9; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_335;
  reg [5:0] depths_10; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_336;
  reg [5:0] depths_11; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_337;
  reg [5:0] depths_12; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_338;
  reg [5:0] depths_13; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_339;
  reg [5:0] depths_14; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_340;
  reg [5:0] depths_15; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_341;
  reg [5:0] depths_16; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_342;
  reg [5:0] depths_17; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_343;
  reg [5:0] depths_18; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_344;
  reg [5:0] depths_19; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_345;
  reg [5:0] depths_20; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_346;
  reg [5:0] depths_21; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_347;
  reg [5:0] depths_22; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_348;
  reg [5:0] depths_23; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_349;
  reg [5:0] depths_24; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_350;
  reg [5:0] depths_25; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_351;
  reg [5:0] depths_26; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_352;
  reg [5:0] depths_27; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_353;
  reg [5:0] depths_28; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_354;
  reg [5:0] depths_29; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_355;
  reg [5:0] depths_30; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_356;
  reg [5:0] depths_31; // @[treeDepthCounter.scala 56:19]
  reg [31:0] _RAND_357;
  reg  state; // @[treeDepthCounter.scala 63:22]
  reg [31:0] _RAND_358;
  wire  _T = ~state; // @[Conditional.scala 37:30]
  wire [6:0] _T_2 = io_inputs_validNodes - 7'h1; // @[treeDepthCounter.scala 82:48]
  wire  _GEN_0 = io_start | state; // @[treeDepthCounter.scala 67:22]
  wire [31:0] _GEN_257 = io_start ? 32'h0 : position; // @[treeDepthCounter.scala 67:22]
  wire [31:0] _GEN_258 = io_start ? 32'h0 : lastNode; // @[treeDepthCounter.scala 67:22]
  wire  _T_4 = charactersVisited >= validCharacters; // @[treeDepthCounter.scala 87:30]
  wire  _T_5 = positionDepth >= lastNodeDepth; // @[treeDepthCounter.scala 91:25]
  wire  _T_6 = positionDepth < lastNodeDepth; // @[treeDepthCounter.scala 91:60]
  wire  _T_7 = ~tpc_io_equal; // @[treeDepthCounter.scala 91:79]
  wire  _T_8 = _T_6 & _T_7; // @[treeDepthCounter.scala 91:76]
  wire  _T_9 = _T_5 | _T_8; // @[treeDepthCounter.scala 91:42]
  wire [8:0] _GEN_265 = 5'h1 == positionDepth[4:0] ? parentNodes_1 : parentNodes_0;
  wire [8:0] _GEN_266 = 5'h2 == positionDepth[4:0] ? parentNodes_2 : _GEN_265;
  wire [8:0] _GEN_267 = 5'h3 == positionDepth[4:0] ? parentNodes_3 : _GEN_266;
  wire [8:0] _GEN_268 = 5'h4 == positionDepth[4:0] ? parentNodes_4 : _GEN_267;
  wire [8:0] _GEN_269 = 5'h5 == positionDepth[4:0] ? parentNodes_5 : _GEN_268;
  wire [8:0] _GEN_270 = 5'h6 == positionDepth[4:0] ? parentNodes_6 : _GEN_269;
  wire [8:0] _GEN_271 = 5'h7 == positionDepth[4:0] ? parentNodes_7 : _GEN_270;
  wire [8:0] _GEN_272 = 5'h8 == positionDepth[4:0] ? parentNodes_8 : _GEN_271;
  wire [8:0] _GEN_273 = 5'h9 == positionDepth[4:0] ? parentNodes_9 : _GEN_272;
  wire [8:0] _GEN_274 = 5'ha == positionDepth[4:0] ? parentNodes_10 : _GEN_273;
  wire [8:0] _GEN_275 = 5'hb == positionDepth[4:0] ? parentNodes_11 : _GEN_274;
  wire [8:0] _GEN_276 = 5'hc == positionDepth[4:0] ? parentNodes_12 : _GEN_275;
  wire [8:0] _GEN_277 = 5'hd == positionDepth[4:0] ? parentNodes_13 : _GEN_276;
  wire [8:0] _GEN_278 = 5'he == positionDepth[4:0] ? parentNodes_14 : _GEN_277;
  wire [8:0] _GEN_279 = 5'hf == positionDepth[4:0] ? parentNodes_15 : _GEN_278;
  wire [8:0] _GEN_280 = 5'h10 == positionDepth[4:0] ? parentNodes_16 : _GEN_279;
  wire [8:0] _GEN_281 = 5'h11 == positionDepth[4:0] ? parentNodes_17 : _GEN_280;
  wire [8:0] _GEN_282 = 5'h12 == positionDepth[4:0] ? parentNodes_18 : _GEN_281;
  wire [8:0] _GEN_283 = 5'h13 == positionDepth[4:0] ? parentNodes_19 : _GEN_282;
  wire [8:0] _GEN_284 = 5'h14 == positionDepth[4:0] ? parentNodes_20 : _GEN_283;
  wire [8:0] _GEN_285 = 5'h15 == positionDepth[4:0] ? parentNodes_21 : _GEN_284;
  wire [8:0] _GEN_286 = 5'h16 == positionDepth[4:0] ? parentNodes_22 : _GEN_285;
  wire [8:0] _GEN_287 = 5'h17 == positionDepth[4:0] ? parentNodes_23 : _GEN_286;
  wire [8:0] _GEN_288 = 5'h18 == positionDepth[4:0] ? parentNodes_24 : _GEN_287;
  wire [8:0] _GEN_289 = 5'h19 == positionDepth[4:0] ? parentNodes_25 : _GEN_288;
  wire [8:0] _GEN_290 = 5'h1a == positionDepth[4:0] ? parentNodes_26 : _GEN_289;
  wire [8:0] _GEN_291 = 5'h1b == positionDepth[4:0] ? parentNodes_27 : _GEN_290;
  wire [8:0] _GEN_292 = 5'h1c == positionDepth[4:0] ? parentNodes_28 : _GEN_291;
  wire [8:0] _GEN_293 = 5'h1d == positionDepth[4:0] ? parentNodes_29 : _GEN_292;
  wire [8:0] _GEN_294 = 5'h1e == positionDepth[4:0] ? parentNodes_30 : _GEN_293;
  wire [8:0] _GEN_295 = 5'h1f == positionDepth[4:0] ? parentNodes_31 : _GEN_294;
  wire  _GEN_297 = 6'h1 == _GEN_295[5:0] ? leftNodeIsCharacter_1 : leftNodeIsCharacter_0; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_298 = 6'h2 == _GEN_295[5:0] ? leftNodeIsCharacter_2 : _GEN_297; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_299 = 6'h3 == _GEN_295[5:0] ? leftNodeIsCharacter_3 : _GEN_298; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_300 = 6'h4 == _GEN_295[5:0] ? leftNodeIsCharacter_4 : _GEN_299; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_301 = 6'h5 == _GEN_295[5:0] ? leftNodeIsCharacter_5 : _GEN_300; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_302 = 6'h6 == _GEN_295[5:0] ? leftNodeIsCharacter_6 : _GEN_301; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_303 = 6'h7 == _GEN_295[5:0] ? leftNodeIsCharacter_7 : _GEN_302; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_304 = 6'h8 == _GEN_295[5:0] ? leftNodeIsCharacter_8 : _GEN_303; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_305 = 6'h9 == _GEN_295[5:0] ? leftNodeIsCharacter_9 : _GEN_304; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_306 = 6'ha == _GEN_295[5:0] ? leftNodeIsCharacter_10 : _GEN_305; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_307 = 6'hb == _GEN_295[5:0] ? leftNodeIsCharacter_11 : _GEN_306; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_308 = 6'hc == _GEN_295[5:0] ? leftNodeIsCharacter_12 : _GEN_307; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_309 = 6'hd == _GEN_295[5:0] ? leftNodeIsCharacter_13 : _GEN_308; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_310 = 6'he == _GEN_295[5:0] ? leftNodeIsCharacter_14 : _GEN_309; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_311 = 6'hf == _GEN_295[5:0] ? leftNodeIsCharacter_15 : _GEN_310; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_312 = 6'h10 == _GEN_295[5:0] ? leftNodeIsCharacter_16 : _GEN_311; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_313 = 6'h11 == _GEN_295[5:0] ? leftNodeIsCharacter_17 : _GEN_312; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_314 = 6'h12 == _GEN_295[5:0] ? leftNodeIsCharacter_18 : _GEN_313; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_315 = 6'h13 == _GEN_295[5:0] ? leftNodeIsCharacter_19 : _GEN_314; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_316 = 6'h14 == _GEN_295[5:0] ? leftNodeIsCharacter_20 : _GEN_315; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_317 = 6'h15 == _GEN_295[5:0] ? leftNodeIsCharacter_21 : _GEN_316; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_318 = 6'h16 == _GEN_295[5:0] ? leftNodeIsCharacter_22 : _GEN_317; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_319 = 6'h17 == _GEN_295[5:0] ? leftNodeIsCharacter_23 : _GEN_318; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_320 = 6'h18 == _GEN_295[5:0] ? leftNodeIsCharacter_24 : _GEN_319; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_321 = 6'h19 == _GEN_295[5:0] ? leftNodeIsCharacter_25 : _GEN_320; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_322 = 6'h1a == _GEN_295[5:0] ? leftNodeIsCharacter_26 : _GEN_321; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_323 = 6'h1b == _GEN_295[5:0] ? leftNodeIsCharacter_27 : _GEN_322; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_324 = 6'h1c == _GEN_295[5:0] ? leftNodeIsCharacter_28 : _GEN_323; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_325 = 6'h1d == _GEN_295[5:0] ? leftNodeIsCharacter_29 : _GEN_324; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_326 = 6'h1e == _GEN_295[5:0] ? leftNodeIsCharacter_30 : _GEN_325; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_327 = 6'h1f == _GEN_295[5:0] ? leftNodeIsCharacter_31 : _GEN_326; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_328 = 6'h20 == _GEN_295[5:0] ? leftNodeIsCharacter_32 : _GEN_327; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_329 = 6'h21 == _GEN_295[5:0] ? leftNodeIsCharacter_33 : _GEN_328; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_330 = 6'h22 == _GEN_295[5:0] ? leftNodeIsCharacter_34 : _GEN_329; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_331 = 6'h23 == _GEN_295[5:0] ? leftNodeIsCharacter_35 : _GEN_330; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_332 = 6'h24 == _GEN_295[5:0] ? leftNodeIsCharacter_36 : _GEN_331; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_333 = 6'h25 == _GEN_295[5:0] ? leftNodeIsCharacter_37 : _GEN_332; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_334 = 6'h26 == _GEN_295[5:0] ? leftNodeIsCharacter_38 : _GEN_333; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_335 = 6'h27 == _GEN_295[5:0] ? leftNodeIsCharacter_39 : _GEN_334; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_336 = 6'h28 == _GEN_295[5:0] ? leftNodeIsCharacter_40 : _GEN_335; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_337 = 6'h29 == _GEN_295[5:0] ? leftNodeIsCharacter_41 : _GEN_336; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_338 = 6'h2a == _GEN_295[5:0] ? leftNodeIsCharacter_42 : _GEN_337; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_339 = 6'h2b == _GEN_295[5:0] ? leftNodeIsCharacter_43 : _GEN_338; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_340 = 6'h2c == _GEN_295[5:0] ? leftNodeIsCharacter_44 : _GEN_339; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_341 = 6'h2d == _GEN_295[5:0] ? leftNodeIsCharacter_45 : _GEN_340; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_342 = 6'h2e == _GEN_295[5:0] ? leftNodeIsCharacter_46 : _GEN_341; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_343 = 6'h2f == _GEN_295[5:0] ? leftNodeIsCharacter_47 : _GEN_342; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_344 = 6'h30 == _GEN_295[5:0] ? leftNodeIsCharacter_48 : _GEN_343; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_345 = 6'h31 == _GEN_295[5:0] ? leftNodeIsCharacter_49 : _GEN_344; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_346 = 6'h32 == _GEN_295[5:0] ? leftNodeIsCharacter_50 : _GEN_345; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_347 = 6'h33 == _GEN_295[5:0] ? leftNodeIsCharacter_51 : _GEN_346; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_348 = 6'h34 == _GEN_295[5:0] ? leftNodeIsCharacter_52 : _GEN_347; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_349 = 6'h35 == _GEN_295[5:0] ? leftNodeIsCharacter_53 : _GEN_348; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_350 = 6'h36 == _GEN_295[5:0] ? leftNodeIsCharacter_54 : _GEN_349; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_351 = 6'h37 == _GEN_295[5:0] ? leftNodeIsCharacter_55 : _GEN_350; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_352 = 6'h38 == _GEN_295[5:0] ? leftNodeIsCharacter_56 : _GEN_351; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_353 = 6'h39 == _GEN_295[5:0] ? leftNodeIsCharacter_57 : _GEN_352; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_354 = 6'h3a == _GEN_295[5:0] ? leftNodeIsCharacter_58 : _GEN_353; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_355 = 6'h3b == _GEN_295[5:0] ? leftNodeIsCharacter_59 : _GEN_354; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_356 = 6'h3c == _GEN_295[5:0] ? leftNodeIsCharacter_60 : _GEN_355; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_357 = 6'h3d == _GEN_295[5:0] ? leftNodeIsCharacter_61 : _GEN_356; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_358 = 6'h3e == _GEN_295[5:0] ? leftNodeIsCharacter_62 : _GEN_357; // @[treeDepthCounter.scala 97:65]
  wire  _GEN_359 = 6'h3f == _GEN_295[5:0] ? leftNodeIsCharacter_63 : _GEN_358; // @[treeDepthCounter.scala 97:65]
  wire [8:0] _GEN_425 = 6'h1 == _GEN_295[5:0] ? leftNode_1 : leftNode_0; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_426 = 6'h2 == _GEN_295[5:0] ? leftNode_2 : _GEN_425; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_427 = 6'h3 == _GEN_295[5:0] ? leftNode_3 : _GEN_426; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_428 = 6'h4 == _GEN_295[5:0] ? leftNode_4 : _GEN_427; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_429 = 6'h5 == _GEN_295[5:0] ? leftNode_5 : _GEN_428; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_430 = 6'h6 == _GEN_295[5:0] ? leftNode_6 : _GEN_429; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_431 = 6'h7 == _GEN_295[5:0] ? leftNode_7 : _GEN_430; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_432 = 6'h8 == _GEN_295[5:0] ? leftNode_8 : _GEN_431; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_433 = 6'h9 == _GEN_295[5:0] ? leftNode_9 : _GEN_432; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_434 = 6'ha == _GEN_295[5:0] ? leftNode_10 : _GEN_433; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_435 = 6'hb == _GEN_295[5:0] ? leftNode_11 : _GEN_434; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_436 = 6'hc == _GEN_295[5:0] ? leftNode_12 : _GEN_435; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_437 = 6'hd == _GEN_295[5:0] ? leftNode_13 : _GEN_436; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_438 = 6'he == _GEN_295[5:0] ? leftNode_14 : _GEN_437; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_439 = 6'hf == _GEN_295[5:0] ? leftNode_15 : _GEN_438; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_440 = 6'h10 == _GEN_295[5:0] ? leftNode_16 : _GEN_439; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_441 = 6'h11 == _GEN_295[5:0] ? leftNode_17 : _GEN_440; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_442 = 6'h12 == _GEN_295[5:0] ? leftNode_18 : _GEN_441; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_443 = 6'h13 == _GEN_295[5:0] ? leftNode_19 : _GEN_442; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_444 = 6'h14 == _GEN_295[5:0] ? leftNode_20 : _GEN_443; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_445 = 6'h15 == _GEN_295[5:0] ? leftNode_21 : _GEN_444; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_446 = 6'h16 == _GEN_295[5:0] ? leftNode_22 : _GEN_445; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_447 = 6'h17 == _GEN_295[5:0] ? leftNode_23 : _GEN_446; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_448 = 6'h18 == _GEN_295[5:0] ? leftNode_24 : _GEN_447; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_449 = 6'h19 == _GEN_295[5:0] ? leftNode_25 : _GEN_448; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_450 = 6'h1a == _GEN_295[5:0] ? leftNode_26 : _GEN_449; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_451 = 6'h1b == _GEN_295[5:0] ? leftNode_27 : _GEN_450; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_452 = 6'h1c == _GEN_295[5:0] ? leftNode_28 : _GEN_451; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_453 = 6'h1d == _GEN_295[5:0] ? leftNode_29 : _GEN_452; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_454 = 6'h1e == _GEN_295[5:0] ? leftNode_30 : _GEN_453; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_455 = 6'h1f == _GEN_295[5:0] ? leftNode_31 : _GEN_454; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_456 = 6'h20 == _GEN_295[5:0] ? leftNode_32 : _GEN_455; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_457 = 6'h21 == _GEN_295[5:0] ? leftNode_33 : _GEN_456; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_458 = 6'h22 == _GEN_295[5:0] ? leftNode_34 : _GEN_457; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_459 = 6'h23 == _GEN_295[5:0] ? leftNode_35 : _GEN_458; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_460 = 6'h24 == _GEN_295[5:0] ? leftNode_36 : _GEN_459; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_461 = 6'h25 == _GEN_295[5:0] ? leftNode_37 : _GEN_460; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_462 = 6'h26 == _GEN_295[5:0] ? leftNode_38 : _GEN_461; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_463 = 6'h27 == _GEN_295[5:0] ? leftNode_39 : _GEN_462; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_464 = 6'h28 == _GEN_295[5:0] ? leftNode_40 : _GEN_463; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_465 = 6'h29 == _GEN_295[5:0] ? leftNode_41 : _GEN_464; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_466 = 6'h2a == _GEN_295[5:0] ? leftNode_42 : _GEN_465; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_467 = 6'h2b == _GEN_295[5:0] ? leftNode_43 : _GEN_466; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_468 = 6'h2c == _GEN_295[5:0] ? leftNode_44 : _GEN_467; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_469 = 6'h2d == _GEN_295[5:0] ? leftNode_45 : _GEN_468; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_470 = 6'h2e == _GEN_295[5:0] ? leftNode_46 : _GEN_469; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_471 = 6'h2f == _GEN_295[5:0] ? leftNode_47 : _GEN_470; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_472 = 6'h30 == _GEN_295[5:0] ? leftNode_48 : _GEN_471; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_473 = 6'h31 == _GEN_295[5:0] ? leftNode_49 : _GEN_472; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_474 = 6'h32 == _GEN_295[5:0] ? leftNode_50 : _GEN_473; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_475 = 6'h33 == _GEN_295[5:0] ? leftNode_51 : _GEN_474; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_476 = 6'h34 == _GEN_295[5:0] ? leftNode_52 : _GEN_475; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_477 = 6'h35 == _GEN_295[5:0] ? leftNode_53 : _GEN_476; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_478 = 6'h36 == _GEN_295[5:0] ? leftNode_54 : _GEN_477; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_479 = 6'h37 == _GEN_295[5:0] ? leftNode_55 : _GEN_478; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_480 = 6'h38 == _GEN_295[5:0] ? leftNode_56 : _GEN_479; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_481 = 6'h39 == _GEN_295[5:0] ? leftNode_57 : _GEN_480; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_482 = 6'h3a == _GEN_295[5:0] ? leftNode_58 : _GEN_481; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_483 = 6'h3b == _GEN_295[5:0] ? leftNode_59 : _GEN_482; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_484 = 6'h3c == _GEN_295[5:0] ? leftNode_60 : _GEN_483; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_485 = 6'h3d == _GEN_295[5:0] ? leftNode_61 : _GEN_484; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_486 = 6'h3e == _GEN_295[5:0] ? leftNode_62 : _GEN_485; // @[treeDepthCounter.scala 99:43]
  wire [8:0] _GEN_487 = 6'h3f == _GEN_295[5:0] ? leftNode_63 : _GEN_486; // @[treeDepthCounter.scala 99:43]
  wire [5:0] _T_17 = positionDepth + 6'h1; // @[treeDepthCounter.scala 102:56]
  wire [5:0] _T_19 = charactersVisited + 6'h1; // @[treeDepthCounter.scala 103:52]
  wire [5:0] _T_23 = 6'h1f - positionDepth; // @[treeDepthCounter.scala 109:82]
  wire [63:0] _T_24 = 64'h1 << _T_23; // @[treeDepthCounter.scala 109:42]
  wire [63:0] _T_25 = ~_T_24; // @[treeDepthCounter.scala 109:36]
  wire [63:0] _GEN_2416 = {{32'd0}, position}; // @[treeDepthCounter.scala 109:34]
  wire [63:0] _T_26 = _GEN_2416 & _T_25; // @[treeDepthCounter.scala 109:34]
  wire  _GEN_553 = 6'h1 == _GEN_295[5:0] ? rightNodeIsCharacter_1 : rightNodeIsCharacter_0; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_554 = 6'h2 == _GEN_295[5:0] ? rightNodeIsCharacter_2 : _GEN_553; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_555 = 6'h3 == _GEN_295[5:0] ? rightNodeIsCharacter_3 : _GEN_554; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_556 = 6'h4 == _GEN_295[5:0] ? rightNodeIsCharacter_4 : _GEN_555; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_557 = 6'h5 == _GEN_295[5:0] ? rightNodeIsCharacter_5 : _GEN_556; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_558 = 6'h6 == _GEN_295[5:0] ? rightNodeIsCharacter_6 : _GEN_557; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_559 = 6'h7 == _GEN_295[5:0] ? rightNodeIsCharacter_7 : _GEN_558; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_560 = 6'h8 == _GEN_295[5:0] ? rightNodeIsCharacter_8 : _GEN_559; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_561 = 6'h9 == _GEN_295[5:0] ? rightNodeIsCharacter_9 : _GEN_560; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_562 = 6'ha == _GEN_295[5:0] ? rightNodeIsCharacter_10 : _GEN_561; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_563 = 6'hb == _GEN_295[5:0] ? rightNodeIsCharacter_11 : _GEN_562; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_564 = 6'hc == _GEN_295[5:0] ? rightNodeIsCharacter_12 : _GEN_563; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_565 = 6'hd == _GEN_295[5:0] ? rightNodeIsCharacter_13 : _GEN_564; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_566 = 6'he == _GEN_295[5:0] ? rightNodeIsCharacter_14 : _GEN_565; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_567 = 6'hf == _GEN_295[5:0] ? rightNodeIsCharacter_15 : _GEN_566; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_568 = 6'h10 == _GEN_295[5:0] ? rightNodeIsCharacter_16 : _GEN_567; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_569 = 6'h11 == _GEN_295[5:0] ? rightNodeIsCharacter_17 : _GEN_568; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_570 = 6'h12 == _GEN_295[5:0] ? rightNodeIsCharacter_18 : _GEN_569; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_571 = 6'h13 == _GEN_295[5:0] ? rightNodeIsCharacter_19 : _GEN_570; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_572 = 6'h14 == _GEN_295[5:0] ? rightNodeIsCharacter_20 : _GEN_571; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_573 = 6'h15 == _GEN_295[5:0] ? rightNodeIsCharacter_21 : _GEN_572; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_574 = 6'h16 == _GEN_295[5:0] ? rightNodeIsCharacter_22 : _GEN_573; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_575 = 6'h17 == _GEN_295[5:0] ? rightNodeIsCharacter_23 : _GEN_574; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_576 = 6'h18 == _GEN_295[5:0] ? rightNodeIsCharacter_24 : _GEN_575; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_577 = 6'h19 == _GEN_295[5:0] ? rightNodeIsCharacter_25 : _GEN_576; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_578 = 6'h1a == _GEN_295[5:0] ? rightNodeIsCharacter_26 : _GEN_577; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_579 = 6'h1b == _GEN_295[5:0] ? rightNodeIsCharacter_27 : _GEN_578; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_580 = 6'h1c == _GEN_295[5:0] ? rightNodeIsCharacter_28 : _GEN_579; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_581 = 6'h1d == _GEN_295[5:0] ? rightNodeIsCharacter_29 : _GEN_580; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_582 = 6'h1e == _GEN_295[5:0] ? rightNodeIsCharacter_30 : _GEN_581; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_583 = 6'h1f == _GEN_295[5:0] ? rightNodeIsCharacter_31 : _GEN_582; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_584 = 6'h20 == _GEN_295[5:0] ? rightNodeIsCharacter_32 : _GEN_583; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_585 = 6'h21 == _GEN_295[5:0] ? rightNodeIsCharacter_33 : _GEN_584; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_586 = 6'h22 == _GEN_295[5:0] ? rightNodeIsCharacter_34 : _GEN_585; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_587 = 6'h23 == _GEN_295[5:0] ? rightNodeIsCharacter_35 : _GEN_586; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_588 = 6'h24 == _GEN_295[5:0] ? rightNodeIsCharacter_36 : _GEN_587; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_589 = 6'h25 == _GEN_295[5:0] ? rightNodeIsCharacter_37 : _GEN_588; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_590 = 6'h26 == _GEN_295[5:0] ? rightNodeIsCharacter_38 : _GEN_589; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_591 = 6'h27 == _GEN_295[5:0] ? rightNodeIsCharacter_39 : _GEN_590; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_592 = 6'h28 == _GEN_295[5:0] ? rightNodeIsCharacter_40 : _GEN_591; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_593 = 6'h29 == _GEN_295[5:0] ? rightNodeIsCharacter_41 : _GEN_592; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_594 = 6'h2a == _GEN_295[5:0] ? rightNodeIsCharacter_42 : _GEN_593; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_595 = 6'h2b == _GEN_295[5:0] ? rightNodeIsCharacter_43 : _GEN_594; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_596 = 6'h2c == _GEN_295[5:0] ? rightNodeIsCharacter_44 : _GEN_595; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_597 = 6'h2d == _GEN_295[5:0] ? rightNodeIsCharacter_45 : _GEN_596; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_598 = 6'h2e == _GEN_295[5:0] ? rightNodeIsCharacter_46 : _GEN_597; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_599 = 6'h2f == _GEN_295[5:0] ? rightNodeIsCharacter_47 : _GEN_598; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_600 = 6'h30 == _GEN_295[5:0] ? rightNodeIsCharacter_48 : _GEN_599; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_601 = 6'h31 == _GEN_295[5:0] ? rightNodeIsCharacter_49 : _GEN_600; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_602 = 6'h32 == _GEN_295[5:0] ? rightNodeIsCharacter_50 : _GEN_601; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_603 = 6'h33 == _GEN_295[5:0] ? rightNodeIsCharacter_51 : _GEN_602; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_604 = 6'h34 == _GEN_295[5:0] ? rightNodeIsCharacter_52 : _GEN_603; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_605 = 6'h35 == _GEN_295[5:0] ? rightNodeIsCharacter_53 : _GEN_604; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_606 = 6'h36 == _GEN_295[5:0] ? rightNodeIsCharacter_54 : _GEN_605; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_607 = 6'h37 == _GEN_295[5:0] ? rightNodeIsCharacter_55 : _GEN_606; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_608 = 6'h38 == _GEN_295[5:0] ? rightNodeIsCharacter_56 : _GEN_607; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_609 = 6'h39 == _GEN_295[5:0] ? rightNodeIsCharacter_57 : _GEN_608; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_610 = 6'h3a == _GEN_295[5:0] ? rightNodeIsCharacter_58 : _GEN_609; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_611 = 6'h3b == _GEN_295[5:0] ? rightNodeIsCharacter_59 : _GEN_610; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_612 = 6'h3c == _GEN_295[5:0] ? rightNodeIsCharacter_60 : _GEN_611; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_613 = 6'h3d == _GEN_295[5:0] ? rightNodeIsCharacter_61 : _GEN_612; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_614 = 6'h3e == _GEN_295[5:0] ? rightNodeIsCharacter_62 : _GEN_613; // @[treeDepthCounter.scala 110:68]
  wire  _GEN_615 = 6'h3f == _GEN_295[5:0] ? rightNodeIsCharacter_63 : _GEN_614; // @[treeDepthCounter.scala 110:68]
  wire [8:0] _GEN_681 = 6'h1 == _GEN_295[5:0] ? rightNode_1 : rightNode_0; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_682 = 6'h2 == _GEN_295[5:0] ? rightNode_2 : _GEN_681; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_683 = 6'h3 == _GEN_295[5:0] ? rightNode_3 : _GEN_682; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_684 = 6'h4 == _GEN_295[5:0] ? rightNode_4 : _GEN_683; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_685 = 6'h5 == _GEN_295[5:0] ? rightNode_5 : _GEN_684; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_686 = 6'h6 == _GEN_295[5:0] ? rightNode_6 : _GEN_685; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_687 = 6'h7 == _GEN_295[5:0] ? rightNode_7 : _GEN_686; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_688 = 6'h8 == _GEN_295[5:0] ? rightNode_8 : _GEN_687; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_689 = 6'h9 == _GEN_295[5:0] ? rightNode_9 : _GEN_688; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_690 = 6'ha == _GEN_295[5:0] ? rightNode_10 : _GEN_689; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_691 = 6'hb == _GEN_295[5:0] ? rightNode_11 : _GEN_690; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_692 = 6'hc == _GEN_295[5:0] ? rightNode_12 : _GEN_691; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_693 = 6'hd == _GEN_295[5:0] ? rightNode_13 : _GEN_692; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_694 = 6'he == _GEN_295[5:0] ? rightNode_14 : _GEN_693; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_695 = 6'hf == _GEN_295[5:0] ? rightNode_15 : _GEN_694; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_696 = 6'h10 == _GEN_295[5:0] ? rightNode_16 : _GEN_695; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_697 = 6'h11 == _GEN_295[5:0] ? rightNode_17 : _GEN_696; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_698 = 6'h12 == _GEN_295[5:0] ? rightNode_18 : _GEN_697; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_699 = 6'h13 == _GEN_295[5:0] ? rightNode_19 : _GEN_698; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_700 = 6'h14 == _GEN_295[5:0] ? rightNode_20 : _GEN_699; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_701 = 6'h15 == _GEN_295[5:0] ? rightNode_21 : _GEN_700; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_702 = 6'h16 == _GEN_295[5:0] ? rightNode_22 : _GEN_701; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_703 = 6'h17 == _GEN_295[5:0] ? rightNode_23 : _GEN_702; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_704 = 6'h18 == _GEN_295[5:0] ? rightNode_24 : _GEN_703; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_705 = 6'h19 == _GEN_295[5:0] ? rightNode_25 : _GEN_704; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_706 = 6'h1a == _GEN_295[5:0] ? rightNode_26 : _GEN_705; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_707 = 6'h1b == _GEN_295[5:0] ? rightNode_27 : _GEN_706; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_708 = 6'h1c == _GEN_295[5:0] ? rightNode_28 : _GEN_707; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_709 = 6'h1d == _GEN_295[5:0] ? rightNode_29 : _GEN_708; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_710 = 6'h1e == _GEN_295[5:0] ? rightNode_30 : _GEN_709; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_711 = 6'h1f == _GEN_295[5:0] ? rightNode_31 : _GEN_710; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_712 = 6'h20 == _GEN_295[5:0] ? rightNode_32 : _GEN_711; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_713 = 6'h21 == _GEN_295[5:0] ? rightNode_33 : _GEN_712; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_714 = 6'h22 == _GEN_295[5:0] ? rightNode_34 : _GEN_713; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_715 = 6'h23 == _GEN_295[5:0] ? rightNode_35 : _GEN_714; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_716 = 6'h24 == _GEN_295[5:0] ? rightNode_36 : _GEN_715; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_717 = 6'h25 == _GEN_295[5:0] ? rightNode_37 : _GEN_716; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_718 = 6'h26 == _GEN_295[5:0] ? rightNode_38 : _GEN_717; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_719 = 6'h27 == _GEN_295[5:0] ? rightNode_39 : _GEN_718; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_720 = 6'h28 == _GEN_295[5:0] ? rightNode_40 : _GEN_719; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_721 = 6'h29 == _GEN_295[5:0] ? rightNode_41 : _GEN_720; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_722 = 6'h2a == _GEN_295[5:0] ? rightNode_42 : _GEN_721; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_723 = 6'h2b == _GEN_295[5:0] ? rightNode_43 : _GEN_722; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_724 = 6'h2c == _GEN_295[5:0] ? rightNode_44 : _GEN_723; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_725 = 6'h2d == _GEN_295[5:0] ? rightNode_45 : _GEN_724; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_726 = 6'h2e == _GEN_295[5:0] ? rightNode_46 : _GEN_725; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_727 = 6'h2f == _GEN_295[5:0] ? rightNode_47 : _GEN_726; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_728 = 6'h30 == _GEN_295[5:0] ? rightNode_48 : _GEN_727; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_729 = 6'h31 == _GEN_295[5:0] ? rightNode_49 : _GEN_728; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_730 = 6'h32 == _GEN_295[5:0] ? rightNode_50 : _GEN_729; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_731 = 6'h33 == _GEN_295[5:0] ? rightNode_51 : _GEN_730; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_732 = 6'h34 == _GEN_295[5:0] ? rightNode_52 : _GEN_731; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_733 = 6'h35 == _GEN_295[5:0] ? rightNode_53 : _GEN_732; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_734 = 6'h36 == _GEN_295[5:0] ? rightNode_54 : _GEN_733; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_735 = 6'h37 == _GEN_295[5:0] ? rightNode_55 : _GEN_734; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_736 = 6'h38 == _GEN_295[5:0] ? rightNode_56 : _GEN_735; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_737 = 6'h39 == _GEN_295[5:0] ? rightNode_57 : _GEN_736; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_738 = 6'h3a == _GEN_295[5:0] ? rightNode_58 : _GEN_737; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_739 = 6'h3b == _GEN_295[5:0] ? rightNode_59 : _GEN_738; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_740 = 6'h3c == _GEN_295[5:0] ? rightNode_60 : _GEN_739; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_741 = 6'h3d == _GEN_295[5:0] ? rightNode_61 : _GEN_740; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_742 = 6'h3e == _GEN_295[5:0] ? rightNode_62 : _GEN_741; // @[treeDepthCounter.scala 113:51]
  wire [8:0] _GEN_743 = 6'h3f == _GEN_295[5:0] ? rightNode_63 : _GEN_742; // @[treeDepthCounter.scala 113:51]
  wire [5:0] _T_40 = charactersVisited + 6'h2; // @[treeDepthCounter.scala 117:54]
  wire [5:0] _T_42 = positionDepth - 6'h1; // @[treeDepthCounter.scala 118:46]
  wire [63:0] _T_46 = _GEN_2416 | _T_24; // @[treeDepthCounter.scala 119:36]
  wire [63:0] _GEN_970 = _GEN_615 ? _T_46 : _T_26; // @[treeDepthCounter.scala 110:68]
  wire [63:0] _GEN_971 = _GEN_615 ? {{32'd0}, position} : _T_46; // @[treeDepthCounter.scala 110:68]
  wire [63:0] _GEN_1198 = _GEN_359 ? _GEN_970 : {{32'd0}, lastNode}; // @[treeDepthCounter.scala 97:65]
  wire [63:0] _GEN_1200 = _GEN_359 ? _GEN_971 : _T_26; // @[treeDepthCounter.scala 97:65]
  wire [31:0] _T_90 = position >> _T_23; // @[treeDepthCounter.scala 153:32]
  wire [31:0] _T_91 = 32'h1 & _T_90; // @[treeDepthCounter.scala 153:20]
  wire  _T_92 = _T_91 == 32'h1; // @[treeDepthCounter.scala 153:91]
  wire [63:0] _GEN_1618 = _T_92 ? {{32'd0}, position} : _T_46; // @[treeDepthCounter.scala 154:15]
  wire [63:0] _GEN_1652 = _GEN_615 ? _T_46 : {{32'd0}, lastNode}; // @[treeDepthCounter.scala 142:66]
  wire [63:0] _GEN_1719 = _GEN_615 ? {{32'd0}, position} : _GEN_1618; // @[treeDepthCounter.scala 142:66]
  wire [63:0] _GEN_1818 = _T_9 ? _GEN_1198 : _GEN_1652; // @[treeDepthCounter.scala 92:11]
  wire [63:0] _GEN_1820 = _T_9 ? _GEN_1200 : _GEN_1719; // @[treeDepthCounter.scala 92:11]
  wire [63:0] _GEN_1920 = _T_4 ? {{32'd0}, lastNode} : _GEN_1818; // @[treeDepthCounter.scala 87:50]
  wire [63:0] _GEN_1922 = _T_4 ? {{32'd0}, position} : _GEN_1820; // @[treeDepthCounter.scala 87:50]
  wire [63:0] _GEN_2022 = state ? _GEN_1920 : {{32'd0}, lastNode}; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_2024 = state ? _GEN_1922 : {{32'd0}, position}; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_2314 = _T ? {{32'd0}, _GEN_257} : _GEN_2024; // @[Conditional.scala 40:58]
  wire [63:0] _GEN_2315 = _T ? {{32'd0}, _GEN_258} : _GEN_2022; // @[Conditional.scala 40:58]
  treePathComparator tpc ( // @[treeDepthCounter.scala 45:19]
    .io_position(tpc_io_position),
    .io_lastNode(tpc_io_lastNode),
    .io_length(tpc_io_length),
    .io_equal(tpc_io_equal)
  );
  assign io_outputs_characters_0 = characters_0; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_1 = characters_1; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_2 = characters_2; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_3 = characters_3; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_4 = characters_4; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_5 = characters_5; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_6 = characters_6; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_7 = characters_7; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_8 = characters_8; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_9 = characters_9; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_10 = characters_10; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_11 = characters_11; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_12 = characters_12; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_13 = characters_13; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_14 = characters_14; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_15 = characters_15; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_16 = characters_16; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_17 = characters_17; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_18 = characters_18; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_19 = characters_19; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_20 = characters_20; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_21 = characters_21; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_22 = characters_22; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_23 = characters_23; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_24 = characters_24; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_25 = characters_25; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_26 = characters_26; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_27 = characters_27; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_28 = characters_28; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_29 = characters_29; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_30 = characters_30; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_characters_31 = characters_31; // @[treeDepthCounter.scala 170:25]
  assign io_outputs_depths_0 = depths_0; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_1 = depths_1; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_2 = depths_2; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_3 = depths_3; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_4 = depths_4; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_5 = depths_5; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_6 = depths_6; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_7 = depths_7; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_8 = depths_8; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_9 = depths_9; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_10 = depths_10; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_11 = depths_11; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_12 = depths_12; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_13 = depths_13; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_14 = depths_14; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_15 = depths_15; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_16 = depths_16; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_17 = depths_17; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_18 = depths_18; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_19 = depths_19; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_20 = depths_20; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_21 = depths_21; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_22 = depths_22; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_23 = depths_23; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_24 = depths_24; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_25 = depths_25; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_26 = depths_26; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_27 = depths_27; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_28 = depths_28; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_29 = depths_29; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_30 = depths_30; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_depths_31 = depths_31; // @[treeDepthCounter.scala 171:21]
  assign io_outputs_validCharacters = validCharacters; // @[treeDepthCounter.scala 172:30]
  assign io_finished = ~state; // @[treeDepthCounter.scala 173:15]
  assign tpc_io_position = position; // @[treeDepthCounter.scala 46:19]
  assign tpc_io_lastNode = lastNode; // @[treeDepthCounter.scala 47:19]
  assign tpc_io_length = positionDepth; // @[treeDepthCounter.scala 48:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  leftNode_0 = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  leftNode_1 = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  leftNode_2 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  leftNode_3 = _RAND_3[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  leftNode_4 = _RAND_4[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  leftNode_5 = _RAND_5[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  leftNode_6 = _RAND_6[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  leftNode_7 = _RAND_7[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  leftNode_8 = _RAND_8[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  leftNode_9 = _RAND_9[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  leftNode_10 = _RAND_10[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  leftNode_11 = _RAND_11[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  leftNode_12 = _RAND_12[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  leftNode_13 = _RAND_13[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  leftNode_14 = _RAND_14[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  leftNode_15 = _RAND_15[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  leftNode_16 = _RAND_16[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  leftNode_17 = _RAND_17[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  leftNode_18 = _RAND_18[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  leftNode_19 = _RAND_19[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  leftNode_20 = _RAND_20[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  leftNode_21 = _RAND_21[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  leftNode_22 = _RAND_22[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  leftNode_23 = _RAND_23[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  leftNode_24 = _RAND_24[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  leftNode_25 = _RAND_25[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  leftNode_26 = _RAND_26[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  leftNode_27 = _RAND_27[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  leftNode_28 = _RAND_28[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  leftNode_29 = _RAND_29[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  leftNode_30 = _RAND_30[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  leftNode_31 = _RAND_31[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  leftNode_32 = _RAND_32[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  leftNode_33 = _RAND_33[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  leftNode_34 = _RAND_34[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  leftNode_35 = _RAND_35[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  leftNode_36 = _RAND_36[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  leftNode_37 = _RAND_37[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  leftNode_38 = _RAND_38[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  leftNode_39 = _RAND_39[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  leftNode_40 = _RAND_40[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  leftNode_41 = _RAND_41[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  leftNode_42 = _RAND_42[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  leftNode_43 = _RAND_43[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  leftNode_44 = _RAND_44[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  leftNode_45 = _RAND_45[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  leftNode_46 = _RAND_46[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  leftNode_47 = _RAND_47[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  leftNode_48 = _RAND_48[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  leftNode_49 = _RAND_49[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  leftNode_50 = _RAND_50[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  leftNode_51 = _RAND_51[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  leftNode_52 = _RAND_52[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  leftNode_53 = _RAND_53[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  leftNode_54 = _RAND_54[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  leftNode_55 = _RAND_55[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  leftNode_56 = _RAND_56[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  leftNode_57 = _RAND_57[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  leftNode_58 = _RAND_58[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  leftNode_59 = _RAND_59[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  leftNode_60 = _RAND_60[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  leftNode_61 = _RAND_61[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  leftNode_62 = _RAND_62[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  leftNode_63 = _RAND_63[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  rightNode_0 = _RAND_64[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  rightNode_1 = _RAND_65[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  rightNode_2 = _RAND_66[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  rightNode_3 = _RAND_67[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  rightNode_4 = _RAND_68[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  rightNode_5 = _RAND_69[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  rightNode_6 = _RAND_70[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  rightNode_7 = _RAND_71[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  rightNode_8 = _RAND_72[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  rightNode_9 = _RAND_73[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  rightNode_10 = _RAND_74[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  rightNode_11 = _RAND_75[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  rightNode_12 = _RAND_76[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  rightNode_13 = _RAND_77[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  rightNode_14 = _RAND_78[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  rightNode_15 = _RAND_79[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  rightNode_16 = _RAND_80[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  rightNode_17 = _RAND_81[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  rightNode_18 = _RAND_82[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  rightNode_19 = _RAND_83[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  rightNode_20 = _RAND_84[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  rightNode_21 = _RAND_85[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  rightNode_22 = _RAND_86[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  rightNode_23 = _RAND_87[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  rightNode_24 = _RAND_88[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  rightNode_25 = _RAND_89[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  rightNode_26 = _RAND_90[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  rightNode_27 = _RAND_91[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  rightNode_28 = _RAND_92[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  rightNode_29 = _RAND_93[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  rightNode_30 = _RAND_94[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  rightNode_31 = _RAND_95[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  rightNode_32 = _RAND_96[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  rightNode_33 = _RAND_97[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  rightNode_34 = _RAND_98[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  rightNode_35 = _RAND_99[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  rightNode_36 = _RAND_100[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  rightNode_37 = _RAND_101[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  rightNode_38 = _RAND_102[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  rightNode_39 = _RAND_103[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  rightNode_40 = _RAND_104[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  rightNode_41 = _RAND_105[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  rightNode_42 = _RAND_106[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  rightNode_43 = _RAND_107[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  rightNode_44 = _RAND_108[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  rightNode_45 = _RAND_109[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  rightNode_46 = _RAND_110[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  rightNode_47 = _RAND_111[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  rightNode_48 = _RAND_112[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  rightNode_49 = _RAND_113[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  rightNode_50 = _RAND_114[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  rightNode_51 = _RAND_115[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  rightNode_52 = _RAND_116[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  rightNode_53 = _RAND_117[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  rightNode_54 = _RAND_118[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  rightNode_55 = _RAND_119[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  rightNode_56 = _RAND_120[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  rightNode_57 = _RAND_121[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  rightNode_58 = _RAND_122[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  rightNode_59 = _RAND_123[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  rightNode_60 = _RAND_124[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  rightNode_61 = _RAND_125[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  rightNode_62 = _RAND_126[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  rightNode_63 = _RAND_127[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  leftNodeIsCharacter_0 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  leftNodeIsCharacter_1 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  leftNodeIsCharacter_2 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  leftNodeIsCharacter_3 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  leftNodeIsCharacter_4 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  leftNodeIsCharacter_5 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  leftNodeIsCharacter_6 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  leftNodeIsCharacter_7 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  leftNodeIsCharacter_8 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  leftNodeIsCharacter_9 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  leftNodeIsCharacter_10 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  leftNodeIsCharacter_11 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  leftNodeIsCharacter_12 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  leftNodeIsCharacter_13 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  leftNodeIsCharacter_14 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  leftNodeIsCharacter_15 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  leftNodeIsCharacter_16 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  leftNodeIsCharacter_17 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  leftNodeIsCharacter_18 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  leftNodeIsCharacter_19 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  leftNodeIsCharacter_20 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  leftNodeIsCharacter_21 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  leftNodeIsCharacter_22 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  leftNodeIsCharacter_23 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  leftNodeIsCharacter_24 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  leftNodeIsCharacter_25 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  leftNodeIsCharacter_26 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  leftNodeIsCharacter_27 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  leftNodeIsCharacter_28 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  leftNodeIsCharacter_29 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  leftNodeIsCharacter_30 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  leftNodeIsCharacter_31 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  leftNodeIsCharacter_32 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  leftNodeIsCharacter_33 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  leftNodeIsCharacter_34 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  leftNodeIsCharacter_35 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  leftNodeIsCharacter_36 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  leftNodeIsCharacter_37 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  leftNodeIsCharacter_38 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  leftNodeIsCharacter_39 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  leftNodeIsCharacter_40 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  leftNodeIsCharacter_41 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  leftNodeIsCharacter_42 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  leftNodeIsCharacter_43 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  leftNodeIsCharacter_44 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  leftNodeIsCharacter_45 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  leftNodeIsCharacter_46 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  leftNodeIsCharacter_47 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  leftNodeIsCharacter_48 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  leftNodeIsCharacter_49 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  leftNodeIsCharacter_50 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  leftNodeIsCharacter_51 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  leftNodeIsCharacter_52 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  leftNodeIsCharacter_53 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  leftNodeIsCharacter_54 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  leftNodeIsCharacter_55 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  leftNodeIsCharacter_56 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  leftNodeIsCharacter_57 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  leftNodeIsCharacter_58 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  leftNodeIsCharacter_59 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  leftNodeIsCharacter_60 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  leftNodeIsCharacter_61 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  leftNodeIsCharacter_62 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  leftNodeIsCharacter_63 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  rightNodeIsCharacter_0 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  rightNodeIsCharacter_1 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  rightNodeIsCharacter_2 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  rightNodeIsCharacter_3 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  rightNodeIsCharacter_4 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  rightNodeIsCharacter_5 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  rightNodeIsCharacter_6 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  rightNodeIsCharacter_7 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  rightNodeIsCharacter_8 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  rightNodeIsCharacter_9 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  rightNodeIsCharacter_10 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  rightNodeIsCharacter_11 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  rightNodeIsCharacter_12 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  rightNodeIsCharacter_13 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  rightNodeIsCharacter_14 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  rightNodeIsCharacter_15 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  rightNodeIsCharacter_16 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  rightNodeIsCharacter_17 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  rightNodeIsCharacter_18 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  rightNodeIsCharacter_19 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  rightNodeIsCharacter_20 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  rightNodeIsCharacter_21 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  rightNodeIsCharacter_22 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  rightNodeIsCharacter_23 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  rightNodeIsCharacter_24 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  rightNodeIsCharacter_25 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  rightNodeIsCharacter_26 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  rightNodeIsCharacter_27 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  rightNodeIsCharacter_28 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  rightNodeIsCharacter_29 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  rightNodeIsCharacter_30 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  rightNodeIsCharacter_31 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  rightNodeIsCharacter_32 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  rightNodeIsCharacter_33 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  rightNodeIsCharacter_34 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  rightNodeIsCharacter_35 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  rightNodeIsCharacter_36 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  rightNodeIsCharacter_37 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  rightNodeIsCharacter_38 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  rightNodeIsCharacter_39 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  rightNodeIsCharacter_40 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  rightNodeIsCharacter_41 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  rightNodeIsCharacter_42 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  rightNodeIsCharacter_43 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  rightNodeIsCharacter_44 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  rightNodeIsCharacter_45 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  rightNodeIsCharacter_46 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  rightNodeIsCharacter_47 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  rightNodeIsCharacter_48 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  rightNodeIsCharacter_49 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  rightNodeIsCharacter_50 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  rightNodeIsCharacter_51 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  rightNodeIsCharacter_52 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  rightNodeIsCharacter_53 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  rightNodeIsCharacter_54 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  rightNodeIsCharacter_55 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  rightNodeIsCharacter_56 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  rightNodeIsCharacter_57 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  rightNodeIsCharacter_58 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  rightNodeIsCharacter_59 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  rightNodeIsCharacter_60 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  rightNodeIsCharacter_61 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  rightNodeIsCharacter_62 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  rightNodeIsCharacter_63 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  validCharacters = _RAND_256[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  charactersVisited = _RAND_257[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  parentNodes_0 = _RAND_258[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  parentNodes_1 = _RAND_259[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  parentNodes_2 = _RAND_260[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  parentNodes_3 = _RAND_261[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  parentNodes_4 = _RAND_262[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  parentNodes_5 = _RAND_263[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  parentNodes_6 = _RAND_264[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  parentNodes_7 = _RAND_265[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  parentNodes_8 = _RAND_266[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  parentNodes_9 = _RAND_267[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  parentNodes_10 = _RAND_268[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  parentNodes_11 = _RAND_269[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  parentNodes_12 = _RAND_270[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  parentNodes_13 = _RAND_271[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  parentNodes_14 = _RAND_272[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  parentNodes_15 = _RAND_273[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  parentNodes_16 = _RAND_274[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  parentNodes_17 = _RAND_275[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  parentNodes_18 = _RAND_276[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  parentNodes_19 = _RAND_277[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  parentNodes_20 = _RAND_278[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  parentNodes_21 = _RAND_279[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  parentNodes_22 = _RAND_280[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  parentNodes_23 = _RAND_281[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  parentNodes_24 = _RAND_282[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  parentNodes_25 = _RAND_283[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  parentNodes_26 = _RAND_284[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  parentNodes_27 = _RAND_285[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  parentNodes_28 = _RAND_286[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  parentNodes_29 = _RAND_287[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  parentNodes_30 = _RAND_288[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  parentNodes_31 = _RAND_289[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  position = _RAND_290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  lastNode = _RAND_291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  positionDepth = _RAND_292[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  lastNodeDepth = _RAND_293[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  characters_0 = _RAND_294[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  characters_1 = _RAND_295[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  characters_2 = _RAND_296[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  characters_3 = _RAND_297[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  characters_4 = _RAND_298[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  characters_5 = _RAND_299[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  characters_6 = _RAND_300[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  characters_7 = _RAND_301[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  characters_8 = _RAND_302[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  characters_9 = _RAND_303[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  characters_10 = _RAND_304[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  characters_11 = _RAND_305[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  characters_12 = _RAND_306[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  characters_13 = _RAND_307[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  characters_14 = _RAND_308[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  characters_15 = _RAND_309[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  characters_16 = _RAND_310[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  characters_17 = _RAND_311[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  characters_18 = _RAND_312[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  characters_19 = _RAND_313[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  characters_20 = _RAND_314[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  characters_21 = _RAND_315[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  characters_22 = _RAND_316[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  characters_23 = _RAND_317[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  characters_24 = _RAND_318[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  characters_25 = _RAND_319[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  characters_26 = _RAND_320[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  characters_27 = _RAND_321[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  characters_28 = _RAND_322[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  characters_29 = _RAND_323[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  characters_30 = _RAND_324[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  characters_31 = _RAND_325[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  depths_0 = _RAND_326[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  depths_1 = _RAND_327[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  depths_2 = _RAND_328[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  depths_3 = _RAND_329[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  depths_4 = _RAND_330[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  depths_5 = _RAND_331[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  depths_6 = _RAND_332[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  depths_7 = _RAND_333[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  depths_8 = _RAND_334[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  depths_9 = _RAND_335[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  depths_10 = _RAND_336[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  depths_11 = _RAND_337[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  depths_12 = _RAND_338[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  depths_13 = _RAND_339[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  depths_14 = _RAND_340[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  depths_15 = _RAND_341[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  depths_16 = _RAND_342[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  depths_17 = _RAND_343[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  depths_18 = _RAND_344[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  depths_19 = _RAND_345[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  depths_20 = _RAND_346[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  depths_21 = _RAND_347[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  depths_22 = _RAND_348[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  depths_23 = _RAND_349[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  depths_24 = _RAND_350[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  depths_25 = _RAND_351[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  depths_26 = _RAND_352[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  depths_27 = _RAND_353[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  depths_28 = _RAND_354[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  depths_29 = _RAND_355[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  depths_30 = _RAND_356[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  depths_31 = _RAND_357[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  state = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T) begin
      if (io_start) begin
        leftNode_0 <= io_inputs_leftNode_0;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_1 <= io_inputs_leftNode_1;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_2 <= io_inputs_leftNode_2;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_3 <= io_inputs_leftNode_3;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_4 <= io_inputs_leftNode_4;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_5 <= io_inputs_leftNode_5;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_6 <= io_inputs_leftNode_6;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_7 <= io_inputs_leftNode_7;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_8 <= io_inputs_leftNode_8;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_9 <= io_inputs_leftNode_9;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_10 <= io_inputs_leftNode_10;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_11 <= io_inputs_leftNode_11;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_12 <= io_inputs_leftNode_12;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_13 <= io_inputs_leftNode_13;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_14 <= io_inputs_leftNode_14;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_15 <= io_inputs_leftNode_15;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_16 <= io_inputs_leftNode_16;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_17 <= io_inputs_leftNode_17;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_18 <= io_inputs_leftNode_18;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_19 <= io_inputs_leftNode_19;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_20 <= io_inputs_leftNode_20;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_21 <= io_inputs_leftNode_21;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_22 <= io_inputs_leftNode_22;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_23 <= io_inputs_leftNode_23;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_24 <= io_inputs_leftNode_24;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_25 <= io_inputs_leftNode_25;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_26 <= io_inputs_leftNode_26;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_27 <= io_inputs_leftNode_27;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_28 <= io_inputs_leftNode_28;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_29 <= io_inputs_leftNode_29;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_30 <= io_inputs_leftNode_30;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_31 <= io_inputs_leftNode_31;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_32 <= io_inputs_leftNode_32;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_33 <= io_inputs_leftNode_33;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_34 <= io_inputs_leftNode_34;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_35 <= io_inputs_leftNode_35;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_36 <= io_inputs_leftNode_36;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_37 <= io_inputs_leftNode_37;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_38 <= io_inputs_leftNode_38;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_39 <= io_inputs_leftNode_39;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_40 <= io_inputs_leftNode_40;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_41 <= io_inputs_leftNode_41;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_42 <= io_inputs_leftNode_42;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_43 <= io_inputs_leftNode_43;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_44 <= io_inputs_leftNode_44;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_45 <= io_inputs_leftNode_45;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_46 <= io_inputs_leftNode_46;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_47 <= io_inputs_leftNode_47;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_48 <= io_inputs_leftNode_48;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_49 <= io_inputs_leftNode_49;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_50 <= io_inputs_leftNode_50;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_51 <= io_inputs_leftNode_51;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_52 <= io_inputs_leftNode_52;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_53 <= io_inputs_leftNode_53;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_54 <= io_inputs_leftNode_54;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_55 <= io_inputs_leftNode_55;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_56 <= io_inputs_leftNode_56;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_57 <= io_inputs_leftNode_57;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_58 <= io_inputs_leftNode_58;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_59 <= io_inputs_leftNode_59;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_60 <= io_inputs_leftNode_60;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_61 <= io_inputs_leftNode_61;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_62 <= io_inputs_leftNode_62;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNode_63 <= io_inputs_leftNode_63;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_0 <= io_inputs_rightNode_0;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_1 <= io_inputs_rightNode_1;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_2 <= io_inputs_rightNode_2;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_3 <= io_inputs_rightNode_3;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_4 <= io_inputs_rightNode_4;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_5 <= io_inputs_rightNode_5;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_6 <= io_inputs_rightNode_6;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_7 <= io_inputs_rightNode_7;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_8 <= io_inputs_rightNode_8;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_9 <= io_inputs_rightNode_9;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_10 <= io_inputs_rightNode_10;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_11 <= io_inputs_rightNode_11;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_12 <= io_inputs_rightNode_12;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_13 <= io_inputs_rightNode_13;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_14 <= io_inputs_rightNode_14;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_15 <= io_inputs_rightNode_15;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_16 <= io_inputs_rightNode_16;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_17 <= io_inputs_rightNode_17;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_18 <= io_inputs_rightNode_18;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_19 <= io_inputs_rightNode_19;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_20 <= io_inputs_rightNode_20;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_21 <= io_inputs_rightNode_21;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_22 <= io_inputs_rightNode_22;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_23 <= io_inputs_rightNode_23;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_24 <= io_inputs_rightNode_24;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_25 <= io_inputs_rightNode_25;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_26 <= io_inputs_rightNode_26;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_27 <= io_inputs_rightNode_27;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_28 <= io_inputs_rightNode_28;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_29 <= io_inputs_rightNode_29;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_30 <= io_inputs_rightNode_30;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_31 <= io_inputs_rightNode_31;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_32 <= io_inputs_rightNode_32;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_33 <= io_inputs_rightNode_33;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_34 <= io_inputs_rightNode_34;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_35 <= io_inputs_rightNode_35;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_36 <= io_inputs_rightNode_36;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_37 <= io_inputs_rightNode_37;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_38 <= io_inputs_rightNode_38;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_39 <= io_inputs_rightNode_39;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_40 <= io_inputs_rightNode_40;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_41 <= io_inputs_rightNode_41;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_42 <= io_inputs_rightNode_42;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_43 <= io_inputs_rightNode_43;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_44 <= io_inputs_rightNode_44;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_45 <= io_inputs_rightNode_45;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_46 <= io_inputs_rightNode_46;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_47 <= io_inputs_rightNode_47;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_48 <= io_inputs_rightNode_48;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_49 <= io_inputs_rightNode_49;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_50 <= io_inputs_rightNode_50;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_51 <= io_inputs_rightNode_51;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_52 <= io_inputs_rightNode_52;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_53 <= io_inputs_rightNode_53;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_54 <= io_inputs_rightNode_54;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_55 <= io_inputs_rightNode_55;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_56 <= io_inputs_rightNode_56;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_57 <= io_inputs_rightNode_57;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_58 <= io_inputs_rightNode_58;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_59 <= io_inputs_rightNode_59;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_60 <= io_inputs_rightNode_60;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_61 <= io_inputs_rightNode_61;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_62 <= io_inputs_rightNode_62;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNode_63 <= io_inputs_rightNode_63;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_0 <= io_inputs_leftNodeIsCharacter_0;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_1 <= io_inputs_leftNodeIsCharacter_1;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_2 <= io_inputs_leftNodeIsCharacter_2;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_3 <= io_inputs_leftNodeIsCharacter_3;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_4 <= io_inputs_leftNodeIsCharacter_4;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_5 <= io_inputs_leftNodeIsCharacter_5;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_6 <= io_inputs_leftNodeIsCharacter_6;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_7 <= io_inputs_leftNodeIsCharacter_7;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_8 <= io_inputs_leftNodeIsCharacter_8;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_9 <= io_inputs_leftNodeIsCharacter_9;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_10 <= io_inputs_leftNodeIsCharacter_10;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_11 <= io_inputs_leftNodeIsCharacter_11;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_12 <= io_inputs_leftNodeIsCharacter_12;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_13 <= io_inputs_leftNodeIsCharacter_13;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_14 <= io_inputs_leftNodeIsCharacter_14;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_15 <= io_inputs_leftNodeIsCharacter_15;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_16 <= io_inputs_leftNodeIsCharacter_16;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_17 <= io_inputs_leftNodeIsCharacter_17;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_18 <= io_inputs_leftNodeIsCharacter_18;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_19 <= io_inputs_leftNodeIsCharacter_19;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_20 <= io_inputs_leftNodeIsCharacter_20;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_21 <= io_inputs_leftNodeIsCharacter_21;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_22 <= io_inputs_leftNodeIsCharacter_22;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_23 <= io_inputs_leftNodeIsCharacter_23;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_24 <= io_inputs_leftNodeIsCharacter_24;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_25 <= io_inputs_leftNodeIsCharacter_25;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_26 <= io_inputs_leftNodeIsCharacter_26;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_27 <= io_inputs_leftNodeIsCharacter_27;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_28 <= io_inputs_leftNodeIsCharacter_28;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_29 <= io_inputs_leftNodeIsCharacter_29;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_30 <= io_inputs_leftNodeIsCharacter_30;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_31 <= io_inputs_leftNodeIsCharacter_31;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_32 <= io_inputs_leftNodeIsCharacter_32;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_33 <= io_inputs_leftNodeIsCharacter_33;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_34 <= io_inputs_leftNodeIsCharacter_34;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_35 <= io_inputs_leftNodeIsCharacter_35;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_36 <= io_inputs_leftNodeIsCharacter_36;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_37 <= io_inputs_leftNodeIsCharacter_37;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_38 <= io_inputs_leftNodeIsCharacter_38;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_39 <= io_inputs_leftNodeIsCharacter_39;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_40 <= io_inputs_leftNodeIsCharacter_40;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_41 <= io_inputs_leftNodeIsCharacter_41;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_42 <= io_inputs_leftNodeIsCharacter_42;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_43 <= io_inputs_leftNodeIsCharacter_43;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_44 <= io_inputs_leftNodeIsCharacter_44;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_45 <= io_inputs_leftNodeIsCharacter_45;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_46 <= io_inputs_leftNodeIsCharacter_46;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_47 <= io_inputs_leftNodeIsCharacter_47;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_48 <= io_inputs_leftNodeIsCharacter_48;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_49 <= io_inputs_leftNodeIsCharacter_49;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_50 <= io_inputs_leftNodeIsCharacter_50;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_51 <= io_inputs_leftNodeIsCharacter_51;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_52 <= io_inputs_leftNodeIsCharacter_52;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_53 <= io_inputs_leftNodeIsCharacter_53;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_54 <= io_inputs_leftNodeIsCharacter_54;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_55 <= io_inputs_leftNodeIsCharacter_55;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_56 <= io_inputs_leftNodeIsCharacter_56;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_57 <= io_inputs_leftNodeIsCharacter_57;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_58 <= io_inputs_leftNodeIsCharacter_58;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_59 <= io_inputs_leftNodeIsCharacter_59;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_60 <= io_inputs_leftNodeIsCharacter_60;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_61 <= io_inputs_leftNodeIsCharacter_61;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_62 <= io_inputs_leftNodeIsCharacter_62;
      end
    end
    if (_T) begin
      if (io_start) begin
        leftNodeIsCharacter_63 <= io_inputs_leftNodeIsCharacter_63;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_0 <= io_inputs_rightNodeIsCharacter_0;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_1 <= io_inputs_rightNodeIsCharacter_1;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_2 <= io_inputs_rightNodeIsCharacter_2;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_3 <= io_inputs_rightNodeIsCharacter_3;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_4 <= io_inputs_rightNodeIsCharacter_4;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_5 <= io_inputs_rightNodeIsCharacter_5;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_6 <= io_inputs_rightNodeIsCharacter_6;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_7 <= io_inputs_rightNodeIsCharacter_7;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_8 <= io_inputs_rightNodeIsCharacter_8;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_9 <= io_inputs_rightNodeIsCharacter_9;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_10 <= io_inputs_rightNodeIsCharacter_10;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_11 <= io_inputs_rightNodeIsCharacter_11;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_12 <= io_inputs_rightNodeIsCharacter_12;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_13 <= io_inputs_rightNodeIsCharacter_13;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_14 <= io_inputs_rightNodeIsCharacter_14;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_15 <= io_inputs_rightNodeIsCharacter_15;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_16 <= io_inputs_rightNodeIsCharacter_16;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_17 <= io_inputs_rightNodeIsCharacter_17;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_18 <= io_inputs_rightNodeIsCharacter_18;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_19 <= io_inputs_rightNodeIsCharacter_19;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_20 <= io_inputs_rightNodeIsCharacter_20;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_21 <= io_inputs_rightNodeIsCharacter_21;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_22 <= io_inputs_rightNodeIsCharacter_22;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_23 <= io_inputs_rightNodeIsCharacter_23;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_24 <= io_inputs_rightNodeIsCharacter_24;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_25 <= io_inputs_rightNodeIsCharacter_25;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_26 <= io_inputs_rightNodeIsCharacter_26;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_27 <= io_inputs_rightNodeIsCharacter_27;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_28 <= io_inputs_rightNodeIsCharacter_28;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_29 <= io_inputs_rightNodeIsCharacter_29;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_30 <= io_inputs_rightNodeIsCharacter_30;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_31 <= io_inputs_rightNodeIsCharacter_31;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_32 <= io_inputs_rightNodeIsCharacter_32;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_33 <= io_inputs_rightNodeIsCharacter_33;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_34 <= io_inputs_rightNodeIsCharacter_34;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_35 <= io_inputs_rightNodeIsCharacter_35;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_36 <= io_inputs_rightNodeIsCharacter_36;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_37 <= io_inputs_rightNodeIsCharacter_37;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_38 <= io_inputs_rightNodeIsCharacter_38;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_39 <= io_inputs_rightNodeIsCharacter_39;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_40 <= io_inputs_rightNodeIsCharacter_40;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_41 <= io_inputs_rightNodeIsCharacter_41;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_42 <= io_inputs_rightNodeIsCharacter_42;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_43 <= io_inputs_rightNodeIsCharacter_43;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_44 <= io_inputs_rightNodeIsCharacter_44;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_45 <= io_inputs_rightNodeIsCharacter_45;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_46 <= io_inputs_rightNodeIsCharacter_46;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_47 <= io_inputs_rightNodeIsCharacter_47;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_48 <= io_inputs_rightNodeIsCharacter_48;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_49 <= io_inputs_rightNodeIsCharacter_49;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_50 <= io_inputs_rightNodeIsCharacter_50;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_51 <= io_inputs_rightNodeIsCharacter_51;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_52 <= io_inputs_rightNodeIsCharacter_52;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_53 <= io_inputs_rightNodeIsCharacter_53;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_54 <= io_inputs_rightNodeIsCharacter_54;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_55 <= io_inputs_rightNodeIsCharacter_55;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_56 <= io_inputs_rightNodeIsCharacter_56;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_57 <= io_inputs_rightNodeIsCharacter_57;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_58 <= io_inputs_rightNodeIsCharacter_58;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_59 <= io_inputs_rightNodeIsCharacter_59;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_60 <= io_inputs_rightNodeIsCharacter_60;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_61 <= io_inputs_rightNodeIsCharacter_61;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_62 <= io_inputs_rightNodeIsCharacter_62;
      end
    end
    if (_T) begin
      if (io_start) begin
        rightNodeIsCharacter_63 <= io_inputs_rightNodeIsCharacter_63;
      end
    end
    if (_T) begin
      if (io_start) begin
        validCharacters <= io_inputs_validCharacters;
      end
    end
    if (_T) begin
      if (io_start) begin
        charactersVisited <= 6'h0;
      end
    end else if (state) begin
      if (!(_T_4)) begin
        if (_T_9) begin
          if (_GEN_359) begin
            if (_GEN_615) begin
              charactersVisited <= _T_40;
            end else begin
              charactersVisited <= _T_19;
            end
          end
        end else if (_GEN_615) begin
          charactersVisited <= _T_19;
        end
      end
    end
    if (_T) begin
      if (io_start) begin
        parentNodes_0 <= {{2'd0}, _T_2};
      end
    end else if (state) begin
      if (!(_T_4)) begin
        if (_T_9) begin
          if (_GEN_359) begin
            if (!(_GEN_615)) begin
              if (5'h0 == _T_17[4:0]) begin
                if (6'h3f == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_63;
                end else if (6'h3e == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_62;
                end else if (6'h3d == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_61;
                end else if (6'h3c == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_60;
                end else if (6'h3b == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_59;
                end else if (6'h3a == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_58;
                end else if (6'h39 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_57;
                end else if (6'h38 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_56;
                end else if (6'h37 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_55;
                end else if (6'h36 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_54;
                end else if (6'h35 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_53;
                end else if (6'h34 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_52;
                end else if (6'h33 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_51;
                end else if (6'h32 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_50;
                end else if (6'h31 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_49;
                end else if (6'h30 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_48;
                end else if (6'h2f == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_47;
                end else if (6'h2e == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_46;
                end else if (6'h2d == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_45;
                end else if (6'h2c == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_44;
                end else if (6'h2b == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_43;
                end else if (6'h2a == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_42;
                end else if (6'h29 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_41;
                end else if (6'h28 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_40;
                end else if (6'h27 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_39;
                end else if (6'h26 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_38;
                end else if (6'h25 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_37;
                end else if (6'h24 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_36;
                end else if (6'h23 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_35;
                end else if (6'h22 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_34;
                end else if (6'h21 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_33;
                end else if (6'h20 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_32;
                end else if (6'h1f == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_31;
                end else if (6'h1e == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_30;
                end else if (6'h1d == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_29;
                end else if (6'h1c == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_28;
                end else if (6'h1b == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_27;
                end else if (6'h1a == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_26;
                end else if (6'h19 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_25;
                end else if (6'h18 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_24;
                end else if (6'h17 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_23;
                end else if (6'h16 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_22;
                end else if (6'h15 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_21;
                end else if (6'h14 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_20;
                end else if (6'h13 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_19;
                end else if (6'h12 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_18;
                end else if (6'h11 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_17;
                end else if (6'h10 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_16;
                end else if (6'hf == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_15;
                end else if (6'he == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_14;
                end else if (6'hd == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_13;
                end else if (6'hc == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_12;
                end else if (6'hb == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_11;
                end else if (6'ha == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_10;
                end else if (6'h9 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_9;
                end else if (6'h8 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_8;
                end else if (6'h7 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_7;
                end else if (6'h6 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_6;
                end else if (6'h5 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_5;
                end else if (6'h4 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_4;
                end else if (6'h3 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_3;
                end else if (6'h2 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_2;
                end else if (6'h1 == _GEN_295[5:0]) begin
                  parentNodes_0 <= rightNode_1;
                end else begin
                  parentNodes_0 <= rightNode_0;
                end
              end
            end
          end else if (5'h0 == _T_17[4:0]) begin
            if (6'h3f == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_63;
            end else if (6'h3e == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_62;
            end else if (6'h3d == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_61;
            end else if (6'h3c == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_60;
            end else if (6'h3b == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_59;
            end else if (6'h3a == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_58;
            end else if (6'h39 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_57;
            end else if (6'h38 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_56;
            end else if (6'h37 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_55;
            end else if (6'h36 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_54;
            end else if (6'h35 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_53;
            end else if (6'h34 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_52;
            end else if (6'h33 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_51;
            end else if (6'h32 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_50;
            end else if (6'h31 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_49;
            end else if (6'h30 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_48;
            end else if (6'h2f == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_47;
            end else if (6'h2e == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_46;
            end else if (6'h2d == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_45;
            end else if (6'h2c == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_44;
            end else if (6'h2b == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_43;
            end else if (6'h2a == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_42;
            end else if (6'h29 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_41;
            end else if (6'h28 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_40;
            end else if (6'h27 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_39;
            end else if (6'h26 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_38;
            end else if (6'h25 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_37;
            end else if (6'h24 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_36;
            end else if (6'h23 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_35;
            end else if (6'h22 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_34;
            end else if (6'h21 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_33;
            end else if (6'h20 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_32;
            end else if (6'h1f == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_31;
            end else if (6'h1e == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_30;
            end else if (6'h1d == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_29;
            end else if (6'h1c == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_28;
            end else if (6'h1b == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_27;
            end else if (6'h1a == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_26;
            end else if (6'h19 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_25;
            end else if (6'h18 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_24;
            end else if (6'h17 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_23;
            end else if (6'h16 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_22;
            end else if (6'h15 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_21;
            end else if (6'h14 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_20;
            end else if (6'h13 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_19;
            end else if (6'h12 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_18;
            end else if (6'h11 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_17;
            end else if (6'h10 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_16;
            end else if (6'hf == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_15;
            end else if (6'he == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_14;
            end else if (6'hd == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_13;
            end else if (6'hc == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_12;
            end else if (6'hb == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_11;
            end else if (6'ha == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_10;
            end else if (6'h9 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_9;
            end else if (6'h8 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_8;
            end else if (6'h7 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_7;
            end else if (6'h6 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_6;
            end else if (6'h5 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_5;
            end else if (6'h4 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_4;
            end else if (6'h3 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_3;
            end else if (6'h2 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_2;
            end else if (6'h1 == _GEN_295[5:0]) begin
              parentNodes_0 <= leftNode_1;
            end else begin
              parentNodes_0 <= leftNode_0;
            end
          end
        end else if (!(_GEN_615)) begin
          if (!(_T_92)) begin
            if (5'h0 == _T_17[4:0]) begin
              if (6'h3f == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_63;
              end else if (6'h3e == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_62;
              end else if (6'h3d == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_61;
              end else if (6'h3c == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_60;
              end else if (6'h3b == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_59;
              end else if (6'h3a == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_58;
              end else if (6'h39 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_57;
              end else if (6'h38 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_56;
              end else if (6'h37 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_55;
              end else if (6'h36 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_54;
              end else if (6'h35 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_53;
              end else if (6'h34 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_52;
              end else if (6'h33 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_51;
              end else if (6'h32 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_50;
              end else if (6'h31 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_49;
              end else if (6'h30 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_48;
              end else if (6'h2f == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_47;
              end else if (6'h2e == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_46;
              end else if (6'h2d == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_45;
              end else if (6'h2c == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_44;
              end else if (6'h2b == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_43;
              end else if (6'h2a == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_42;
              end else if (6'h29 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_41;
              end else if (6'h28 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_40;
              end else if (6'h27 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_39;
              end else if (6'h26 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_38;
              end else if (6'h25 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_37;
              end else if (6'h24 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_36;
              end else if (6'h23 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_35;
              end else if (6'h22 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_34;
              end else if (6'h21 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_33;
              end else if (6'h20 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_32;
              end else if (6'h1f == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_31;
              end else if (6'h1e == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_30;
              end else if (6'h1d == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_29;
              end else if (6'h1c == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_28;
              end else if (6'h1b == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_27;
              end else if (6'h1a == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_26;
              end else if (6'h19 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_25;
              end else if (6'h18 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_24;
              end else if (6'h17 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_23;
              end else if (6'h16 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_22;
              end else if (6'h15 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_21;
              end else if (6'h14 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_20;
              end else if (6'h13 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_19;
              end else if (6'h12 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_18;
              end else if (6'h11 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_17;
              end else if (6'h10 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_16;
              end else if (6'hf == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_15;
              end else if (6'he == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_14;
              end else if (6'hd == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_13;
              end else if (6'hc == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_12;
              end else if (6'hb == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_11;
              end else if (6'ha == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_10;
              end else if (6'h9 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_9;
              end else if (6'h8 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_8;
              end else if (6'h7 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_7;
              end else if (6'h6 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_6;
              end else if (6'h5 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_5;
              end else if (6'h4 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_4;
              end else if (6'h3 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_3;
              end else if (6'h2 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_2;
              end else if (6'h1 == _GEN_295[5:0]) begin
                parentNodes_0 <= rightNode_1;
              end else begin
                parentNodes_0 <= rightNode_0;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h1 == _T_17[4:0]) begin
                  if (6'h3f == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_63;
                  end else if (6'h3e == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_62;
                  end else if (6'h3d == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_61;
                  end else if (6'h3c == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_60;
                  end else if (6'h3b == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_59;
                  end else if (6'h3a == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_58;
                  end else if (6'h39 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_57;
                  end else if (6'h38 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_56;
                  end else if (6'h37 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_55;
                  end else if (6'h36 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_54;
                  end else if (6'h35 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_53;
                  end else if (6'h34 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_52;
                  end else if (6'h33 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_51;
                  end else if (6'h32 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_50;
                  end else if (6'h31 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_49;
                  end else if (6'h30 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_48;
                  end else if (6'h2f == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_47;
                  end else if (6'h2e == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_46;
                  end else if (6'h2d == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_45;
                  end else if (6'h2c == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_44;
                  end else if (6'h2b == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_43;
                  end else if (6'h2a == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_42;
                  end else if (6'h29 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_41;
                  end else if (6'h28 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_40;
                  end else if (6'h27 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_39;
                  end else if (6'h26 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_38;
                  end else if (6'h25 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_37;
                  end else if (6'h24 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_36;
                  end else if (6'h23 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_35;
                  end else if (6'h22 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_34;
                  end else if (6'h21 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_33;
                  end else if (6'h20 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_32;
                  end else if (6'h1f == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_31;
                  end else if (6'h1e == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_30;
                  end else if (6'h1d == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_29;
                  end else if (6'h1c == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_28;
                  end else if (6'h1b == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_27;
                  end else if (6'h1a == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_26;
                  end else if (6'h19 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_25;
                  end else if (6'h18 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_24;
                  end else if (6'h17 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_23;
                  end else if (6'h16 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_22;
                  end else if (6'h15 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_21;
                  end else if (6'h14 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_20;
                  end else if (6'h13 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_19;
                  end else if (6'h12 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_18;
                  end else if (6'h11 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_17;
                  end else if (6'h10 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_16;
                  end else if (6'hf == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_15;
                  end else if (6'he == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_14;
                  end else if (6'hd == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_13;
                  end else if (6'hc == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_12;
                  end else if (6'hb == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_11;
                  end else if (6'ha == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_10;
                  end else if (6'h9 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_9;
                  end else if (6'h8 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_8;
                  end else if (6'h7 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_7;
                  end else if (6'h6 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_6;
                  end else if (6'h5 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_5;
                  end else if (6'h4 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_4;
                  end else if (6'h3 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_3;
                  end else if (6'h2 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_2;
                  end else if (6'h1 == _GEN_295[5:0]) begin
                    parentNodes_1 <= rightNode_1;
                  end else begin
                    parentNodes_1 <= rightNode_0;
                  end
                end
              end
            end else if (5'h1 == _T_17[4:0]) begin
              if (6'h3f == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_63;
              end else if (6'h3e == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_62;
              end else if (6'h3d == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_61;
              end else if (6'h3c == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_60;
              end else if (6'h3b == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_59;
              end else if (6'h3a == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_58;
              end else if (6'h39 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_57;
              end else if (6'h38 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_56;
              end else if (6'h37 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_55;
              end else if (6'h36 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_54;
              end else if (6'h35 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_53;
              end else if (6'h34 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_52;
              end else if (6'h33 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_51;
              end else if (6'h32 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_50;
              end else if (6'h31 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_49;
              end else if (6'h30 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_48;
              end else if (6'h2f == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_47;
              end else if (6'h2e == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_46;
              end else if (6'h2d == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_45;
              end else if (6'h2c == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_44;
              end else if (6'h2b == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_43;
              end else if (6'h2a == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_42;
              end else if (6'h29 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_41;
              end else if (6'h28 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_40;
              end else if (6'h27 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_39;
              end else if (6'h26 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_38;
              end else if (6'h25 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_37;
              end else if (6'h24 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_36;
              end else if (6'h23 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_35;
              end else if (6'h22 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_34;
              end else if (6'h21 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_33;
              end else if (6'h20 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_32;
              end else if (6'h1f == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_31;
              end else if (6'h1e == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_30;
              end else if (6'h1d == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_29;
              end else if (6'h1c == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_28;
              end else if (6'h1b == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_27;
              end else if (6'h1a == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_26;
              end else if (6'h19 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_25;
              end else if (6'h18 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_24;
              end else if (6'h17 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_23;
              end else if (6'h16 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_22;
              end else if (6'h15 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_21;
              end else if (6'h14 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_20;
              end else if (6'h13 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_19;
              end else if (6'h12 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_18;
              end else if (6'h11 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_17;
              end else if (6'h10 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_16;
              end else if (6'hf == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_15;
              end else if (6'he == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_14;
              end else if (6'hd == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_13;
              end else if (6'hc == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_12;
              end else if (6'hb == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_11;
              end else if (6'ha == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_10;
              end else if (6'h9 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_9;
              end else if (6'h8 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_8;
              end else if (6'h7 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_7;
              end else if (6'h6 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_6;
              end else if (6'h5 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_5;
              end else if (6'h4 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_4;
              end else if (6'h3 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_3;
              end else if (6'h2 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_2;
              end else if (6'h1 == _GEN_295[5:0]) begin
                parentNodes_1 <= leftNode_1;
              end else begin
                parentNodes_1 <= leftNode_0;
              end
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h1 == _T_17[4:0]) begin
                if (6'h3f == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_63;
                end else if (6'h3e == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_62;
                end else if (6'h3d == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_61;
                end else if (6'h3c == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_60;
                end else if (6'h3b == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_59;
                end else if (6'h3a == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_58;
                end else if (6'h39 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_57;
                end else if (6'h38 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_56;
                end else if (6'h37 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_55;
                end else if (6'h36 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_54;
                end else if (6'h35 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_53;
                end else if (6'h34 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_52;
                end else if (6'h33 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_51;
                end else if (6'h32 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_50;
                end else if (6'h31 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_49;
                end else if (6'h30 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_48;
                end else if (6'h2f == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_47;
                end else if (6'h2e == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_46;
                end else if (6'h2d == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_45;
                end else if (6'h2c == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_44;
                end else if (6'h2b == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_43;
                end else if (6'h2a == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_42;
                end else if (6'h29 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_41;
                end else if (6'h28 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_40;
                end else if (6'h27 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_39;
                end else if (6'h26 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_38;
                end else if (6'h25 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_37;
                end else if (6'h24 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_36;
                end else if (6'h23 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_35;
                end else if (6'h22 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_34;
                end else if (6'h21 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_33;
                end else if (6'h20 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_32;
                end else if (6'h1f == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_31;
                end else if (6'h1e == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_30;
                end else if (6'h1d == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_29;
                end else if (6'h1c == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_28;
                end else if (6'h1b == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_27;
                end else if (6'h1a == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_26;
                end else if (6'h19 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_25;
                end else if (6'h18 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_24;
                end else if (6'h17 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_23;
                end else if (6'h16 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_22;
                end else if (6'h15 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_21;
                end else if (6'h14 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_20;
                end else if (6'h13 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_19;
                end else if (6'h12 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_18;
                end else if (6'h11 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_17;
                end else if (6'h10 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_16;
                end else if (6'hf == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_15;
                end else if (6'he == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_14;
                end else if (6'hd == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_13;
                end else if (6'hc == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_12;
                end else if (6'hb == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_11;
                end else if (6'ha == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_10;
                end else if (6'h9 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_9;
                end else if (6'h8 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_8;
                end else if (6'h7 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_7;
                end else if (6'h6 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_6;
                end else if (6'h5 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_5;
                end else if (6'h4 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_4;
                end else if (6'h3 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_3;
                end else if (6'h2 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_2;
                end else if (6'h1 == _GEN_295[5:0]) begin
                  parentNodes_1 <= rightNode_1;
                end else begin
                  parentNodes_1 <= rightNode_0;
                end
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h2 == _T_17[4:0]) begin
                  parentNodes_2 <= _GEN_743;
                end
              end
            end else if (5'h2 == _T_17[4:0]) begin
              if (6'h3f == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_63;
              end else if (6'h3e == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_62;
              end else if (6'h3d == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_61;
              end else if (6'h3c == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_60;
              end else if (6'h3b == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_59;
              end else if (6'h3a == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_58;
              end else if (6'h39 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_57;
              end else if (6'h38 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_56;
              end else if (6'h37 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_55;
              end else if (6'h36 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_54;
              end else if (6'h35 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_53;
              end else if (6'h34 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_52;
              end else if (6'h33 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_51;
              end else if (6'h32 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_50;
              end else if (6'h31 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_49;
              end else if (6'h30 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_48;
              end else if (6'h2f == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_47;
              end else if (6'h2e == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_46;
              end else if (6'h2d == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_45;
              end else if (6'h2c == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_44;
              end else if (6'h2b == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_43;
              end else if (6'h2a == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_42;
              end else if (6'h29 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_41;
              end else if (6'h28 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_40;
              end else if (6'h27 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_39;
              end else if (6'h26 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_38;
              end else if (6'h25 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_37;
              end else if (6'h24 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_36;
              end else if (6'h23 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_35;
              end else if (6'h22 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_34;
              end else if (6'h21 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_33;
              end else if (6'h20 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_32;
              end else if (6'h1f == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_31;
              end else if (6'h1e == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_30;
              end else if (6'h1d == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_29;
              end else if (6'h1c == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_28;
              end else if (6'h1b == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_27;
              end else if (6'h1a == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_26;
              end else if (6'h19 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_25;
              end else if (6'h18 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_24;
              end else if (6'h17 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_23;
              end else if (6'h16 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_22;
              end else if (6'h15 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_21;
              end else if (6'h14 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_20;
              end else if (6'h13 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_19;
              end else if (6'h12 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_18;
              end else if (6'h11 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_17;
              end else if (6'h10 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_16;
              end else if (6'hf == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_15;
              end else if (6'he == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_14;
              end else if (6'hd == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_13;
              end else if (6'hc == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_12;
              end else if (6'hb == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_11;
              end else if (6'ha == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_10;
              end else if (6'h9 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_9;
              end else if (6'h8 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_8;
              end else if (6'h7 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_7;
              end else if (6'h6 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_6;
              end else if (6'h5 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_5;
              end else if (6'h4 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_4;
              end else if (6'h3 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_3;
              end else if (6'h2 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_2;
              end else if (6'h1 == _GEN_295[5:0]) begin
                parentNodes_2 <= leftNode_1;
              end else begin
                parentNodes_2 <= leftNode_0;
              end
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h2 == _T_17[4:0]) begin
                parentNodes_2 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h3 == _T_17[4:0]) begin
                  parentNodes_3 <= _GEN_743;
                end
              end
            end else if (5'h3 == _T_17[4:0]) begin
              if (6'h3f == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_63;
              end else if (6'h3e == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_62;
              end else if (6'h3d == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_61;
              end else if (6'h3c == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_60;
              end else if (6'h3b == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_59;
              end else if (6'h3a == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_58;
              end else if (6'h39 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_57;
              end else if (6'h38 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_56;
              end else if (6'h37 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_55;
              end else if (6'h36 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_54;
              end else if (6'h35 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_53;
              end else if (6'h34 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_52;
              end else if (6'h33 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_51;
              end else if (6'h32 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_50;
              end else if (6'h31 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_49;
              end else if (6'h30 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_48;
              end else if (6'h2f == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_47;
              end else if (6'h2e == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_46;
              end else if (6'h2d == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_45;
              end else if (6'h2c == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_44;
              end else if (6'h2b == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_43;
              end else if (6'h2a == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_42;
              end else if (6'h29 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_41;
              end else if (6'h28 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_40;
              end else if (6'h27 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_39;
              end else if (6'h26 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_38;
              end else if (6'h25 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_37;
              end else if (6'h24 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_36;
              end else if (6'h23 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_35;
              end else if (6'h22 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_34;
              end else if (6'h21 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_33;
              end else if (6'h20 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_32;
              end else if (6'h1f == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_31;
              end else if (6'h1e == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_30;
              end else if (6'h1d == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_29;
              end else if (6'h1c == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_28;
              end else if (6'h1b == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_27;
              end else if (6'h1a == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_26;
              end else if (6'h19 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_25;
              end else if (6'h18 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_24;
              end else if (6'h17 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_23;
              end else if (6'h16 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_22;
              end else if (6'h15 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_21;
              end else if (6'h14 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_20;
              end else if (6'h13 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_19;
              end else if (6'h12 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_18;
              end else if (6'h11 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_17;
              end else if (6'h10 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_16;
              end else if (6'hf == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_15;
              end else if (6'he == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_14;
              end else if (6'hd == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_13;
              end else if (6'hc == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_12;
              end else if (6'hb == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_11;
              end else if (6'ha == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_10;
              end else if (6'h9 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_9;
              end else if (6'h8 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_8;
              end else if (6'h7 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_7;
              end else if (6'h6 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_6;
              end else if (6'h5 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_5;
              end else if (6'h4 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_4;
              end else if (6'h3 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_3;
              end else if (6'h2 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_2;
              end else if (6'h1 == _GEN_295[5:0]) begin
                parentNodes_3 <= leftNode_1;
              end else begin
                parentNodes_3 <= leftNode_0;
              end
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h3 == _T_17[4:0]) begin
                parentNodes_3 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h4 == _T_17[4:0]) begin
                  parentNodes_4 <= _GEN_743;
                end
              end
            end else if (5'h4 == _T_17[4:0]) begin
              parentNodes_4 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h4 == _T_17[4:0]) begin
                parentNodes_4 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h5 == _T_17[4:0]) begin
                  parentNodes_5 <= _GEN_743;
                end
              end
            end else if (5'h5 == _T_17[4:0]) begin
              parentNodes_5 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h5 == _T_17[4:0]) begin
                parentNodes_5 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h6 == _T_17[4:0]) begin
                  parentNodes_6 <= _GEN_743;
                end
              end
            end else if (5'h6 == _T_17[4:0]) begin
              parentNodes_6 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h6 == _T_17[4:0]) begin
                parentNodes_6 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h7 == _T_17[4:0]) begin
                  parentNodes_7 <= _GEN_743;
                end
              end
            end else if (5'h7 == _T_17[4:0]) begin
              parentNodes_7 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h7 == _T_17[4:0]) begin
                parentNodes_7 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h8 == _T_17[4:0]) begin
                  parentNodes_8 <= _GEN_743;
                end
              end
            end else if (5'h8 == _T_17[4:0]) begin
              parentNodes_8 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h8 == _T_17[4:0]) begin
                parentNodes_8 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h9 == _T_17[4:0]) begin
                  parentNodes_9 <= _GEN_743;
                end
              end
            end else if (5'h9 == _T_17[4:0]) begin
              parentNodes_9 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h9 == _T_17[4:0]) begin
                parentNodes_9 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'ha == _T_17[4:0]) begin
                  parentNodes_10 <= _GEN_743;
                end
              end
            end else if (5'ha == _T_17[4:0]) begin
              parentNodes_10 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'ha == _T_17[4:0]) begin
                parentNodes_10 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'hb == _T_17[4:0]) begin
                  parentNodes_11 <= _GEN_743;
                end
              end
            end else if (5'hb == _T_17[4:0]) begin
              parentNodes_11 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'hb == _T_17[4:0]) begin
                parentNodes_11 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'hc == _T_17[4:0]) begin
                  parentNodes_12 <= _GEN_743;
                end
              end
            end else if (5'hc == _T_17[4:0]) begin
              parentNodes_12 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'hc == _T_17[4:0]) begin
                parentNodes_12 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'hd == _T_17[4:0]) begin
                  parentNodes_13 <= _GEN_743;
                end
              end
            end else if (5'hd == _T_17[4:0]) begin
              parentNodes_13 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'hd == _T_17[4:0]) begin
                parentNodes_13 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'he == _T_17[4:0]) begin
                  parentNodes_14 <= _GEN_743;
                end
              end
            end else if (5'he == _T_17[4:0]) begin
              parentNodes_14 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'he == _T_17[4:0]) begin
                parentNodes_14 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'hf == _T_17[4:0]) begin
                  parentNodes_15 <= _GEN_743;
                end
              end
            end else if (5'hf == _T_17[4:0]) begin
              parentNodes_15 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'hf == _T_17[4:0]) begin
                parentNodes_15 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h10 == _T_17[4:0]) begin
                  parentNodes_16 <= _GEN_743;
                end
              end
            end else if (5'h10 == _T_17[4:0]) begin
              parentNodes_16 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h10 == _T_17[4:0]) begin
                parentNodes_16 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h11 == _T_17[4:0]) begin
                  parentNodes_17 <= _GEN_743;
                end
              end
            end else if (5'h11 == _T_17[4:0]) begin
              parentNodes_17 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h11 == _T_17[4:0]) begin
                parentNodes_17 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h12 == _T_17[4:0]) begin
                  parentNodes_18 <= _GEN_743;
                end
              end
            end else if (5'h12 == _T_17[4:0]) begin
              parentNodes_18 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h12 == _T_17[4:0]) begin
                parentNodes_18 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h13 == _T_17[4:0]) begin
                  parentNodes_19 <= _GEN_743;
                end
              end
            end else if (5'h13 == _T_17[4:0]) begin
              parentNodes_19 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h13 == _T_17[4:0]) begin
                parentNodes_19 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h14 == _T_17[4:0]) begin
                  parentNodes_20 <= _GEN_743;
                end
              end
            end else if (5'h14 == _T_17[4:0]) begin
              parentNodes_20 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h14 == _T_17[4:0]) begin
                parentNodes_20 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h15 == _T_17[4:0]) begin
                  parentNodes_21 <= _GEN_743;
                end
              end
            end else if (5'h15 == _T_17[4:0]) begin
              parentNodes_21 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h15 == _T_17[4:0]) begin
                parentNodes_21 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h16 == _T_17[4:0]) begin
                  parentNodes_22 <= _GEN_743;
                end
              end
            end else if (5'h16 == _T_17[4:0]) begin
              parentNodes_22 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h16 == _T_17[4:0]) begin
                parentNodes_22 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h17 == _T_17[4:0]) begin
                  parentNodes_23 <= _GEN_743;
                end
              end
            end else if (5'h17 == _T_17[4:0]) begin
              parentNodes_23 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h17 == _T_17[4:0]) begin
                parentNodes_23 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h18 == _T_17[4:0]) begin
                  parentNodes_24 <= _GEN_743;
                end
              end
            end else if (5'h18 == _T_17[4:0]) begin
              parentNodes_24 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h18 == _T_17[4:0]) begin
                parentNodes_24 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h19 == _T_17[4:0]) begin
                  parentNodes_25 <= _GEN_743;
                end
              end
            end else if (5'h19 == _T_17[4:0]) begin
              parentNodes_25 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h19 == _T_17[4:0]) begin
                parentNodes_25 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h1a == _T_17[4:0]) begin
                  parentNodes_26 <= _GEN_743;
                end
              end
            end else if (5'h1a == _T_17[4:0]) begin
              parentNodes_26 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h1a == _T_17[4:0]) begin
                parentNodes_26 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h1b == _T_17[4:0]) begin
                  parentNodes_27 <= _GEN_743;
                end
              end
            end else if (5'h1b == _T_17[4:0]) begin
              parentNodes_27 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h1b == _T_17[4:0]) begin
                parentNodes_27 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h1c == _T_17[4:0]) begin
                  parentNodes_28 <= _GEN_743;
                end
              end
            end else if (5'h1c == _T_17[4:0]) begin
              parentNodes_28 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h1c == _T_17[4:0]) begin
                parentNodes_28 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h1d == _T_17[4:0]) begin
                  parentNodes_29 <= _GEN_743;
                end
              end
            end else if (5'h1d == _T_17[4:0]) begin
              parentNodes_29 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h1d == _T_17[4:0]) begin
                parentNodes_29 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h1e == _T_17[4:0]) begin
                  parentNodes_30 <= _GEN_743;
                end
              end
            end else if (5'h1e == _T_17[4:0]) begin
              parentNodes_30 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h1e == _T_17[4:0]) begin
                parentNodes_30 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (!(_GEN_615)) begin
                if (5'h1f == _T_17[4:0]) begin
                  parentNodes_31 <= _GEN_743;
                end
              end
            end else if (5'h1f == _T_17[4:0]) begin
              parentNodes_31 <= _GEN_487;
            end
          end else if (!(_GEN_615)) begin
            if (!(_T_92)) begin
              if (5'h1f == _T_17[4:0]) begin
                parentNodes_31 <= _GEN_743;
              end
            end
          end
        end
      end
    end
    position <= _GEN_2314[31:0];
    lastNode <= _GEN_2315[31:0];
    if (_T) begin
      if (io_start) begin
        positionDepth <= 6'h0;
      end
    end else if (state) begin
      if (!(_T_4)) begin
        if (_T_9) begin
          if (_GEN_359) begin
            if (_GEN_615) begin
              positionDepth <= _T_42;
            end else begin
              positionDepth <= _T_17;
            end
          end else begin
            positionDepth <= _T_17;
          end
        end else if (_GEN_615) begin
          positionDepth <= _T_42;
        end else if (_T_92) begin
          positionDepth <= _T_42;
        end else begin
          positionDepth <= _T_17;
        end
      end
    end
    if (_T) begin
      if (io_start) begin
        lastNodeDepth <= 6'h0;
      end
    end else if (state) begin
      if (!(_T_4)) begin
        if (_T_9) begin
          if (_GEN_359) begin
            lastNodeDepth <= _T_17;
          end
        end else if (_GEN_615) begin
          lastNodeDepth <= _T_17;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h0 == _T_19[4:0]) begin
                  characters_0 <= _GEN_743;
                end else if (5'h0 == charactersVisited[4:0]) begin
                  characters_0 <= _GEN_487;
                end
              end else if (5'h0 == charactersVisited[4:0]) begin
                characters_0 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h0 == charactersVisited[4:0]) begin
              characters_0 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h1 == _T_19[4:0]) begin
                  characters_1 <= _GEN_743;
                end else if (5'h1 == charactersVisited[4:0]) begin
                  characters_1 <= _GEN_487;
                end
              end else if (5'h1 == charactersVisited[4:0]) begin
                characters_1 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h1 == charactersVisited[4:0]) begin
              characters_1 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h2 == _T_19[4:0]) begin
                  characters_2 <= _GEN_743;
                end else if (5'h2 == charactersVisited[4:0]) begin
                  characters_2 <= _GEN_487;
                end
              end else if (5'h2 == charactersVisited[4:0]) begin
                characters_2 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h2 == charactersVisited[4:0]) begin
              characters_2 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h3 == _T_19[4:0]) begin
                  characters_3 <= _GEN_743;
                end else if (5'h3 == charactersVisited[4:0]) begin
                  characters_3 <= _GEN_487;
                end
              end else if (5'h3 == charactersVisited[4:0]) begin
                characters_3 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h3 == charactersVisited[4:0]) begin
              characters_3 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h4 == _T_19[4:0]) begin
                  characters_4 <= _GEN_743;
                end else if (5'h4 == charactersVisited[4:0]) begin
                  characters_4 <= _GEN_487;
                end
              end else if (5'h4 == charactersVisited[4:0]) begin
                characters_4 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h4 == charactersVisited[4:0]) begin
              characters_4 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h5 == _T_19[4:0]) begin
                  characters_5 <= _GEN_743;
                end else if (5'h5 == charactersVisited[4:0]) begin
                  characters_5 <= _GEN_487;
                end
              end else if (5'h5 == charactersVisited[4:0]) begin
                characters_5 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h5 == charactersVisited[4:0]) begin
              characters_5 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h6 == _T_19[4:0]) begin
                  characters_6 <= _GEN_743;
                end else if (5'h6 == charactersVisited[4:0]) begin
                  characters_6 <= _GEN_487;
                end
              end else if (5'h6 == charactersVisited[4:0]) begin
                characters_6 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h6 == charactersVisited[4:0]) begin
              characters_6 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h7 == _T_19[4:0]) begin
                  characters_7 <= _GEN_743;
                end else if (5'h7 == charactersVisited[4:0]) begin
                  characters_7 <= _GEN_487;
                end
              end else if (5'h7 == charactersVisited[4:0]) begin
                characters_7 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h7 == charactersVisited[4:0]) begin
              characters_7 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h8 == _T_19[4:0]) begin
                  characters_8 <= _GEN_743;
                end else if (5'h8 == charactersVisited[4:0]) begin
                  characters_8 <= _GEN_487;
                end
              end else if (5'h8 == charactersVisited[4:0]) begin
                characters_8 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h8 == charactersVisited[4:0]) begin
              characters_8 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h9 == _T_19[4:0]) begin
                  characters_9 <= _GEN_743;
                end else if (5'h9 == charactersVisited[4:0]) begin
                  characters_9 <= _GEN_487;
                end
              end else if (5'h9 == charactersVisited[4:0]) begin
                characters_9 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h9 == charactersVisited[4:0]) begin
              characters_9 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'ha == _T_19[4:0]) begin
                  characters_10 <= _GEN_743;
                end else if (5'ha == charactersVisited[4:0]) begin
                  characters_10 <= _GEN_487;
                end
              end else if (5'ha == charactersVisited[4:0]) begin
                characters_10 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'ha == charactersVisited[4:0]) begin
              characters_10 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'hb == _T_19[4:0]) begin
                  characters_11 <= _GEN_743;
                end else if (5'hb == charactersVisited[4:0]) begin
                  characters_11 <= _GEN_487;
                end
              end else if (5'hb == charactersVisited[4:0]) begin
                characters_11 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'hb == charactersVisited[4:0]) begin
              characters_11 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'hc == _T_19[4:0]) begin
                  characters_12 <= _GEN_743;
                end else if (5'hc == charactersVisited[4:0]) begin
                  characters_12 <= _GEN_487;
                end
              end else if (5'hc == charactersVisited[4:0]) begin
                characters_12 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'hc == charactersVisited[4:0]) begin
              characters_12 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'hd == _T_19[4:0]) begin
                  characters_13 <= _GEN_743;
                end else if (5'hd == charactersVisited[4:0]) begin
                  characters_13 <= _GEN_487;
                end
              end else if (5'hd == charactersVisited[4:0]) begin
                characters_13 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'hd == charactersVisited[4:0]) begin
              characters_13 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'he == _T_19[4:0]) begin
                  characters_14 <= _GEN_743;
                end else if (5'he == charactersVisited[4:0]) begin
                  characters_14 <= _GEN_487;
                end
              end else if (5'he == charactersVisited[4:0]) begin
                characters_14 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'he == charactersVisited[4:0]) begin
              characters_14 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'hf == _T_19[4:0]) begin
                  characters_15 <= _GEN_743;
                end else if (5'hf == charactersVisited[4:0]) begin
                  characters_15 <= _GEN_487;
                end
              end else if (5'hf == charactersVisited[4:0]) begin
                characters_15 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'hf == charactersVisited[4:0]) begin
              characters_15 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h10 == _T_19[4:0]) begin
                  characters_16 <= _GEN_743;
                end else if (5'h10 == charactersVisited[4:0]) begin
                  characters_16 <= _GEN_487;
                end
              end else if (5'h10 == charactersVisited[4:0]) begin
                characters_16 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h10 == charactersVisited[4:0]) begin
              characters_16 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h11 == _T_19[4:0]) begin
                  characters_17 <= _GEN_743;
                end else if (5'h11 == charactersVisited[4:0]) begin
                  characters_17 <= _GEN_487;
                end
              end else if (5'h11 == charactersVisited[4:0]) begin
                characters_17 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h11 == charactersVisited[4:0]) begin
              characters_17 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h12 == _T_19[4:0]) begin
                  characters_18 <= _GEN_743;
                end else if (5'h12 == charactersVisited[4:0]) begin
                  characters_18 <= _GEN_487;
                end
              end else if (5'h12 == charactersVisited[4:0]) begin
                characters_18 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h12 == charactersVisited[4:0]) begin
              characters_18 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h13 == _T_19[4:0]) begin
                  characters_19 <= _GEN_743;
                end else if (5'h13 == charactersVisited[4:0]) begin
                  characters_19 <= _GEN_487;
                end
              end else if (5'h13 == charactersVisited[4:0]) begin
                characters_19 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h13 == charactersVisited[4:0]) begin
              characters_19 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h14 == _T_19[4:0]) begin
                  characters_20 <= _GEN_743;
                end else if (5'h14 == charactersVisited[4:0]) begin
                  characters_20 <= _GEN_487;
                end
              end else if (5'h14 == charactersVisited[4:0]) begin
                characters_20 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h14 == charactersVisited[4:0]) begin
              characters_20 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h15 == _T_19[4:0]) begin
                  characters_21 <= _GEN_743;
                end else if (5'h15 == charactersVisited[4:0]) begin
                  characters_21 <= _GEN_487;
                end
              end else if (5'h15 == charactersVisited[4:0]) begin
                characters_21 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h15 == charactersVisited[4:0]) begin
              characters_21 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h16 == _T_19[4:0]) begin
                  characters_22 <= _GEN_743;
                end else if (5'h16 == charactersVisited[4:0]) begin
                  characters_22 <= _GEN_487;
                end
              end else if (5'h16 == charactersVisited[4:0]) begin
                characters_22 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h16 == charactersVisited[4:0]) begin
              characters_22 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h17 == _T_19[4:0]) begin
                  characters_23 <= _GEN_743;
                end else if (5'h17 == charactersVisited[4:0]) begin
                  characters_23 <= _GEN_487;
                end
              end else if (5'h17 == charactersVisited[4:0]) begin
                characters_23 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h17 == charactersVisited[4:0]) begin
              characters_23 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h18 == _T_19[4:0]) begin
                  characters_24 <= _GEN_743;
                end else if (5'h18 == charactersVisited[4:0]) begin
                  characters_24 <= _GEN_487;
                end
              end else if (5'h18 == charactersVisited[4:0]) begin
                characters_24 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h18 == charactersVisited[4:0]) begin
              characters_24 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h19 == _T_19[4:0]) begin
                  characters_25 <= _GEN_743;
                end else if (5'h19 == charactersVisited[4:0]) begin
                  characters_25 <= _GEN_487;
                end
              end else if (5'h19 == charactersVisited[4:0]) begin
                characters_25 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h19 == charactersVisited[4:0]) begin
              characters_25 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h1a == _T_19[4:0]) begin
                  characters_26 <= _GEN_743;
                end else if (5'h1a == charactersVisited[4:0]) begin
                  characters_26 <= _GEN_487;
                end
              end else if (5'h1a == charactersVisited[4:0]) begin
                characters_26 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h1a == charactersVisited[4:0]) begin
              characters_26 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h1b == _T_19[4:0]) begin
                  characters_27 <= _GEN_743;
                end else if (5'h1b == charactersVisited[4:0]) begin
                  characters_27 <= _GEN_487;
                end
              end else if (5'h1b == charactersVisited[4:0]) begin
                characters_27 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h1b == charactersVisited[4:0]) begin
              characters_27 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h1c == _T_19[4:0]) begin
                  characters_28 <= _GEN_743;
                end else if (5'h1c == charactersVisited[4:0]) begin
                  characters_28 <= _GEN_487;
                end
              end else if (5'h1c == charactersVisited[4:0]) begin
                characters_28 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h1c == charactersVisited[4:0]) begin
              characters_28 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h1d == _T_19[4:0]) begin
                  characters_29 <= _GEN_743;
                end else if (5'h1d == charactersVisited[4:0]) begin
                  characters_29 <= _GEN_487;
                end
              end else if (5'h1d == charactersVisited[4:0]) begin
                characters_29 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h1d == charactersVisited[4:0]) begin
              characters_29 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h1e == _T_19[4:0]) begin
                  characters_30 <= _GEN_743;
                end else if (5'h1e == charactersVisited[4:0]) begin
                  characters_30 <= _GEN_487;
                end
              end else if (5'h1e == charactersVisited[4:0]) begin
                characters_30 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h1e == charactersVisited[4:0]) begin
              characters_30 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h1f == _T_19[4:0]) begin
                  characters_31 <= _GEN_743;
                end else if (5'h1f == charactersVisited[4:0]) begin
                  characters_31 <= _GEN_487;
                end
              end else if (5'h1f == charactersVisited[4:0]) begin
                characters_31 <= _GEN_487;
              end
            end
          end else if (_GEN_615) begin
            if (5'h1f == charactersVisited[4:0]) begin
              characters_31 <= _GEN_743;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h0 == _T_19[4:0]) begin
                  depths_0 <= _T_17;
                end else if (5'h0 == charactersVisited[4:0]) begin
                  depths_0 <= _T_17;
                end
              end else if (5'h0 == charactersVisited[4:0]) begin
                depths_0 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h0 == charactersVisited[4:0]) begin
              depths_0 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h1 == _T_19[4:0]) begin
                  depths_1 <= _T_17;
                end else if (5'h1 == charactersVisited[4:0]) begin
                  depths_1 <= _T_17;
                end
              end else if (5'h1 == charactersVisited[4:0]) begin
                depths_1 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h1 == charactersVisited[4:0]) begin
              depths_1 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h2 == _T_19[4:0]) begin
                  depths_2 <= _T_17;
                end else if (5'h2 == charactersVisited[4:0]) begin
                  depths_2 <= _T_17;
                end
              end else if (5'h2 == charactersVisited[4:0]) begin
                depths_2 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h2 == charactersVisited[4:0]) begin
              depths_2 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h3 == _T_19[4:0]) begin
                  depths_3 <= _T_17;
                end else if (5'h3 == charactersVisited[4:0]) begin
                  depths_3 <= _T_17;
                end
              end else if (5'h3 == charactersVisited[4:0]) begin
                depths_3 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h3 == charactersVisited[4:0]) begin
              depths_3 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h4 == _T_19[4:0]) begin
                  depths_4 <= _T_17;
                end else if (5'h4 == charactersVisited[4:0]) begin
                  depths_4 <= _T_17;
                end
              end else if (5'h4 == charactersVisited[4:0]) begin
                depths_4 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h4 == charactersVisited[4:0]) begin
              depths_4 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h5 == _T_19[4:0]) begin
                  depths_5 <= _T_17;
                end else if (5'h5 == charactersVisited[4:0]) begin
                  depths_5 <= _T_17;
                end
              end else if (5'h5 == charactersVisited[4:0]) begin
                depths_5 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h5 == charactersVisited[4:0]) begin
              depths_5 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h6 == _T_19[4:0]) begin
                  depths_6 <= _T_17;
                end else if (5'h6 == charactersVisited[4:0]) begin
                  depths_6 <= _T_17;
                end
              end else if (5'h6 == charactersVisited[4:0]) begin
                depths_6 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h6 == charactersVisited[4:0]) begin
              depths_6 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h7 == _T_19[4:0]) begin
                  depths_7 <= _T_17;
                end else if (5'h7 == charactersVisited[4:0]) begin
                  depths_7 <= _T_17;
                end
              end else if (5'h7 == charactersVisited[4:0]) begin
                depths_7 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h7 == charactersVisited[4:0]) begin
              depths_7 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h8 == _T_19[4:0]) begin
                  depths_8 <= _T_17;
                end else if (5'h8 == charactersVisited[4:0]) begin
                  depths_8 <= _T_17;
                end
              end else if (5'h8 == charactersVisited[4:0]) begin
                depths_8 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h8 == charactersVisited[4:0]) begin
              depths_8 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h9 == _T_19[4:0]) begin
                  depths_9 <= _T_17;
                end else if (5'h9 == charactersVisited[4:0]) begin
                  depths_9 <= _T_17;
                end
              end else if (5'h9 == charactersVisited[4:0]) begin
                depths_9 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h9 == charactersVisited[4:0]) begin
              depths_9 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'ha == _T_19[4:0]) begin
                  depths_10 <= _T_17;
                end else if (5'ha == charactersVisited[4:0]) begin
                  depths_10 <= _T_17;
                end
              end else if (5'ha == charactersVisited[4:0]) begin
                depths_10 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'ha == charactersVisited[4:0]) begin
              depths_10 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'hb == _T_19[4:0]) begin
                  depths_11 <= _T_17;
                end else if (5'hb == charactersVisited[4:0]) begin
                  depths_11 <= _T_17;
                end
              end else if (5'hb == charactersVisited[4:0]) begin
                depths_11 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'hb == charactersVisited[4:0]) begin
              depths_11 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'hc == _T_19[4:0]) begin
                  depths_12 <= _T_17;
                end else if (5'hc == charactersVisited[4:0]) begin
                  depths_12 <= _T_17;
                end
              end else if (5'hc == charactersVisited[4:0]) begin
                depths_12 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'hc == charactersVisited[4:0]) begin
              depths_12 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'hd == _T_19[4:0]) begin
                  depths_13 <= _T_17;
                end else if (5'hd == charactersVisited[4:0]) begin
                  depths_13 <= _T_17;
                end
              end else if (5'hd == charactersVisited[4:0]) begin
                depths_13 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'hd == charactersVisited[4:0]) begin
              depths_13 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'he == _T_19[4:0]) begin
                  depths_14 <= _T_17;
                end else if (5'he == charactersVisited[4:0]) begin
                  depths_14 <= _T_17;
                end
              end else if (5'he == charactersVisited[4:0]) begin
                depths_14 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'he == charactersVisited[4:0]) begin
              depths_14 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'hf == _T_19[4:0]) begin
                  depths_15 <= _T_17;
                end else if (5'hf == charactersVisited[4:0]) begin
                  depths_15 <= _T_17;
                end
              end else if (5'hf == charactersVisited[4:0]) begin
                depths_15 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'hf == charactersVisited[4:0]) begin
              depths_15 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h10 == _T_19[4:0]) begin
                  depths_16 <= _T_17;
                end else if (5'h10 == charactersVisited[4:0]) begin
                  depths_16 <= _T_17;
                end
              end else if (5'h10 == charactersVisited[4:0]) begin
                depths_16 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h10 == charactersVisited[4:0]) begin
              depths_16 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h11 == _T_19[4:0]) begin
                  depths_17 <= _T_17;
                end else if (5'h11 == charactersVisited[4:0]) begin
                  depths_17 <= _T_17;
                end
              end else if (5'h11 == charactersVisited[4:0]) begin
                depths_17 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h11 == charactersVisited[4:0]) begin
              depths_17 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h12 == _T_19[4:0]) begin
                  depths_18 <= _T_17;
                end else if (5'h12 == charactersVisited[4:0]) begin
                  depths_18 <= _T_17;
                end
              end else if (5'h12 == charactersVisited[4:0]) begin
                depths_18 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h12 == charactersVisited[4:0]) begin
              depths_18 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h13 == _T_19[4:0]) begin
                  depths_19 <= _T_17;
                end else if (5'h13 == charactersVisited[4:0]) begin
                  depths_19 <= _T_17;
                end
              end else if (5'h13 == charactersVisited[4:0]) begin
                depths_19 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h13 == charactersVisited[4:0]) begin
              depths_19 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h14 == _T_19[4:0]) begin
                  depths_20 <= _T_17;
                end else if (5'h14 == charactersVisited[4:0]) begin
                  depths_20 <= _T_17;
                end
              end else if (5'h14 == charactersVisited[4:0]) begin
                depths_20 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h14 == charactersVisited[4:0]) begin
              depths_20 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h15 == _T_19[4:0]) begin
                  depths_21 <= _T_17;
                end else if (5'h15 == charactersVisited[4:0]) begin
                  depths_21 <= _T_17;
                end
              end else if (5'h15 == charactersVisited[4:0]) begin
                depths_21 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h15 == charactersVisited[4:0]) begin
              depths_21 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h16 == _T_19[4:0]) begin
                  depths_22 <= _T_17;
                end else if (5'h16 == charactersVisited[4:0]) begin
                  depths_22 <= _T_17;
                end
              end else if (5'h16 == charactersVisited[4:0]) begin
                depths_22 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h16 == charactersVisited[4:0]) begin
              depths_22 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h17 == _T_19[4:0]) begin
                  depths_23 <= _T_17;
                end else if (5'h17 == charactersVisited[4:0]) begin
                  depths_23 <= _T_17;
                end
              end else if (5'h17 == charactersVisited[4:0]) begin
                depths_23 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h17 == charactersVisited[4:0]) begin
              depths_23 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h18 == _T_19[4:0]) begin
                  depths_24 <= _T_17;
                end else if (5'h18 == charactersVisited[4:0]) begin
                  depths_24 <= _T_17;
                end
              end else if (5'h18 == charactersVisited[4:0]) begin
                depths_24 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h18 == charactersVisited[4:0]) begin
              depths_24 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h19 == _T_19[4:0]) begin
                  depths_25 <= _T_17;
                end else if (5'h19 == charactersVisited[4:0]) begin
                  depths_25 <= _T_17;
                end
              end else if (5'h19 == charactersVisited[4:0]) begin
                depths_25 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h19 == charactersVisited[4:0]) begin
              depths_25 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h1a == _T_19[4:0]) begin
                  depths_26 <= _T_17;
                end else if (5'h1a == charactersVisited[4:0]) begin
                  depths_26 <= _T_17;
                end
              end else if (5'h1a == charactersVisited[4:0]) begin
                depths_26 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h1a == charactersVisited[4:0]) begin
              depths_26 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h1b == _T_19[4:0]) begin
                  depths_27 <= _T_17;
                end else if (5'h1b == charactersVisited[4:0]) begin
                  depths_27 <= _T_17;
                end
              end else if (5'h1b == charactersVisited[4:0]) begin
                depths_27 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h1b == charactersVisited[4:0]) begin
              depths_27 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h1c == _T_19[4:0]) begin
                  depths_28 <= _T_17;
                end else if (5'h1c == charactersVisited[4:0]) begin
                  depths_28 <= _T_17;
                end
              end else if (5'h1c == charactersVisited[4:0]) begin
                depths_28 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h1c == charactersVisited[4:0]) begin
              depths_28 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h1d == _T_19[4:0]) begin
                  depths_29 <= _T_17;
                end else if (5'h1d == charactersVisited[4:0]) begin
                  depths_29 <= _T_17;
                end
              end else if (5'h1d == charactersVisited[4:0]) begin
                depths_29 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h1d == charactersVisited[4:0]) begin
              depths_29 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h1e == _T_19[4:0]) begin
                  depths_30 <= _T_17;
                end else if (5'h1e == charactersVisited[4:0]) begin
                  depths_30 <= _T_17;
                end
              end else if (5'h1e == charactersVisited[4:0]) begin
                depths_30 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h1e == charactersVisited[4:0]) begin
              depths_30 <= _T_17;
            end
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (!(_T_4)) begin
          if (_T_9) begin
            if (_GEN_359) begin
              if (_GEN_615) begin
                if (5'h1f == _T_19[4:0]) begin
                  depths_31 <= _T_17;
                end else if (5'h1f == charactersVisited[4:0]) begin
                  depths_31 <= _T_17;
                end
              end else if (5'h1f == charactersVisited[4:0]) begin
                depths_31 <= _T_17;
              end
            end
          end else if (_GEN_615) begin
            if (5'h1f == charactersVisited[4:0]) begin
              depths_31 <= _T_17;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T) begin
      state <= _GEN_0;
    end else if (state) begin
      if (_T_4) begin
        state <= 1'h0;
      end
    end
  end
endmodule
module sort(
  input        clock,
  input        reset,
  input        io_start,
  input  [8:0] io_inputs_characters_0,
  input  [8:0] io_inputs_characters_1,
  input  [8:0] io_inputs_characters_2,
  input  [8:0] io_inputs_characters_3,
  input  [8:0] io_inputs_characters_4,
  input  [8:0] io_inputs_characters_5,
  input  [8:0] io_inputs_characters_6,
  input  [8:0] io_inputs_characters_7,
  input  [8:0] io_inputs_characters_8,
  input  [8:0] io_inputs_characters_9,
  input  [8:0] io_inputs_characters_10,
  input  [8:0] io_inputs_characters_11,
  input  [8:0] io_inputs_characters_12,
  input  [8:0] io_inputs_characters_13,
  input  [8:0] io_inputs_characters_14,
  input  [8:0] io_inputs_characters_15,
  input  [8:0] io_inputs_characters_16,
  input  [8:0] io_inputs_characters_17,
  input  [8:0] io_inputs_characters_18,
  input  [8:0] io_inputs_characters_19,
  input  [8:0] io_inputs_characters_20,
  input  [8:0] io_inputs_characters_21,
  input  [8:0] io_inputs_characters_22,
  input  [8:0] io_inputs_characters_23,
  input  [8:0] io_inputs_characters_24,
  input  [8:0] io_inputs_characters_25,
  input  [8:0] io_inputs_characters_26,
  input  [8:0] io_inputs_characters_27,
  input  [8:0] io_inputs_characters_28,
  input  [8:0] io_inputs_characters_29,
  input  [8:0] io_inputs_characters_30,
  input  [8:0] io_inputs_characters_31,
  input  [5:0] io_inputs_depths_0,
  input  [5:0] io_inputs_depths_1,
  input  [5:0] io_inputs_depths_2,
  input  [5:0] io_inputs_depths_3,
  input  [5:0] io_inputs_depths_4,
  input  [5:0] io_inputs_depths_5,
  input  [5:0] io_inputs_depths_6,
  input  [5:0] io_inputs_depths_7,
  input  [5:0] io_inputs_depths_8,
  input  [5:0] io_inputs_depths_9,
  input  [5:0] io_inputs_depths_10,
  input  [5:0] io_inputs_depths_11,
  input  [5:0] io_inputs_depths_12,
  input  [5:0] io_inputs_depths_13,
  input  [5:0] io_inputs_depths_14,
  input  [5:0] io_inputs_depths_15,
  input  [5:0] io_inputs_depths_16,
  input  [5:0] io_inputs_depths_17,
  input  [5:0] io_inputs_depths_18,
  input  [5:0] io_inputs_depths_19,
  input  [5:0] io_inputs_depths_20,
  input  [5:0] io_inputs_depths_21,
  input  [5:0] io_inputs_depths_22,
  input  [5:0] io_inputs_depths_23,
  input  [5:0] io_inputs_depths_24,
  input  [5:0] io_inputs_depths_25,
  input  [5:0] io_inputs_depths_26,
  input  [5:0] io_inputs_depths_27,
  input  [5:0] io_inputs_depths_28,
  input  [5:0] io_inputs_depths_29,
  input  [5:0] io_inputs_depths_30,
  input  [5:0] io_inputs_depths_31,
  input  [5:0] io_inputs_validCharacters,
  output [7:0] io_outputs_outputData_0,
  output [7:0] io_outputs_outputData_1,
  output [7:0] io_outputs_outputData_2,
  output [7:0] io_outputs_outputData_3,
  output [7:0] io_outputs_outputData_4,
  output [7:0] io_outputs_outputData_5,
  output [7:0] io_outputs_outputData_6,
  output [7:0] io_outputs_outputData_7,
  output [7:0] io_outputs_outputData_8,
  output [7:0] io_outputs_outputData_9,
  output [7:0] io_outputs_outputData_10,
  output [7:0] io_outputs_outputData_11,
  output [7:0] io_outputs_outputData_12,
  output [7:0] io_outputs_outputData_13,
  output [7:0] io_outputs_outputData_14,
  output [7:0] io_outputs_outputData_15,
  output [7:0] io_outputs_outputData_16,
  output [7:0] io_outputs_outputData_17,
  output [7:0] io_outputs_outputData_18,
  output [7:0] io_outputs_outputData_19,
  output [7:0] io_outputs_outputData_20,
  output [7:0] io_outputs_outputData_21,
  output [7:0] io_outputs_outputData_22,
  output [7:0] io_outputs_outputData_23,
  output [7:0] io_outputs_outputData_24,
  output [7:0] io_outputs_outputData_25,
  output [7:0] io_outputs_outputData_26,
  output [7:0] io_outputs_outputData_27,
  output [7:0] io_outputs_outputData_28,
  output [7:0] io_outputs_outputData_29,
  output [7:0] io_outputs_outputData_30,
  output [7:0] io_outputs_outputData_31,
  output [8:0] io_outputs_outputTags_0,
  output [8:0] io_outputs_outputTags_1,
  output [8:0] io_outputs_outputTags_2,
  output [8:0] io_outputs_outputTags_3,
  output [8:0] io_outputs_outputTags_4,
  output [8:0] io_outputs_outputTags_5,
  output [8:0] io_outputs_outputTags_6,
  output [8:0] io_outputs_outputTags_7,
  output [8:0] io_outputs_outputTags_8,
  output [8:0] io_outputs_outputTags_9,
  output [8:0] io_outputs_outputTags_10,
  output [8:0] io_outputs_outputTags_11,
  output [8:0] io_outputs_outputTags_12,
  output [8:0] io_outputs_outputTags_13,
  output [8:0] io_outputs_outputTags_14,
  output [8:0] io_outputs_outputTags_15,
  output [8:0] io_outputs_outputTags_16,
  output [8:0] io_outputs_outputTags_17,
  output [8:0] io_outputs_outputTags_18,
  output [8:0] io_outputs_outputTags_19,
  output [8:0] io_outputs_outputTags_20,
  output [8:0] io_outputs_outputTags_21,
  output [8:0] io_outputs_outputTags_22,
  output [8:0] io_outputs_outputTags_23,
  output [8:0] io_outputs_outputTags_24,
  output [8:0] io_outputs_outputTags_25,
  output [8:0] io_outputs_outputTags_26,
  output [8:0] io_outputs_outputTags_27,
  output [8:0] io_outputs_outputTags_28,
  output [8:0] io_outputs_outputTags_29,
  output [8:0] io_outputs_outputTags_30,
  output [8:0] io_outputs_outputTags_31,
  output [5:0] io_outputs_itemNumber,
  output       io_finished
);
  reg  state; // @[sort.scala 25:22]
  reg [31:0] _RAND_0;
  reg [5:0] iteration; // @[sort.scala 27:22]
  reg [31:0] _RAND_1;
  reg [8:0] sortData_0; // @[sort.scala 28:21]
  reg [31:0] _RAND_2;
  reg [8:0] sortData_1; // @[sort.scala 28:21]
  reg [31:0] _RAND_3;
  reg [8:0] sortData_2; // @[sort.scala 28:21]
  reg [31:0] _RAND_4;
  reg [8:0] sortData_3; // @[sort.scala 28:21]
  reg [31:0] _RAND_5;
  reg [8:0] sortData_4; // @[sort.scala 28:21]
  reg [31:0] _RAND_6;
  reg [8:0] sortData_5; // @[sort.scala 28:21]
  reg [31:0] _RAND_7;
  reg [8:0] sortData_6; // @[sort.scala 28:21]
  reg [31:0] _RAND_8;
  reg [8:0] sortData_7; // @[sort.scala 28:21]
  reg [31:0] _RAND_9;
  reg [8:0] sortData_8; // @[sort.scala 28:21]
  reg [31:0] _RAND_10;
  reg [8:0] sortData_9; // @[sort.scala 28:21]
  reg [31:0] _RAND_11;
  reg [8:0] sortData_10; // @[sort.scala 28:21]
  reg [31:0] _RAND_12;
  reg [8:0] sortData_11; // @[sort.scala 28:21]
  reg [31:0] _RAND_13;
  reg [8:0] sortData_12; // @[sort.scala 28:21]
  reg [31:0] _RAND_14;
  reg [8:0] sortData_13; // @[sort.scala 28:21]
  reg [31:0] _RAND_15;
  reg [8:0] sortData_14; // @[sort.scala 28:21]
  reg [31:0] _RAND_16;
  reg [8:0] sortData_15; // @[sort.scala 28:21]
  reg [31:0] _RAND_17;
  reg [8:0] sortData_16; // @[sort.scala 28:21]
  reg [31:0] _RAND_18;
  reg [8:0] sortData_17; // @[sort.scala 28:21]
  reg [31:0] _RAND_19;
  reg [8:0] sortData_18; // @[sort.scala 28:21]
  reg [31:0] _RAND_20;
  reg [8:0] sortData_19; // @[sort.scala 28:21]
  reg [31:0] _RAND_21;
  reg [8:0] sortData_20; // @[sort.scala 28:21]
  reg [31:0] _RAND_22;
  reg [8:0] sortData_21; // @[sort.scala 28:21]
  reg [31:0] _RAND_23;
  reg [8:0] sortData_22; // @[sort.scala 28:21]
  reg [31:0] _RAND_24;
  reg [8:0] sortData_23; // @[sort.scala 28:21]
  reg [31:0] _RAND_25;
  reg [8:0] sortData_24; // @[sort.scala 28:21]
  reg [31:0] _RAND_26;
  reg [8:0] sortData_25; // @[sort.scala 28:21]
  reg [31:0] _RAND_27;
  reg [8:0] sortData_26; // @[sort.scala 28:21]
  reg [31:0] _RAND_28;
  reg [8:0] sortData_27; // @[sort.scala 28:21]
  reg [31:0] _RAND_29;
  reg [8:0] sortData_28; // @[sort.scala 28:21]
  reg [31:0] _RAND_30;
  reg [8:0] sortData_29; // @[sort.scala 28:21]
  reg [31:0] _RAND_31;
  reg [8:0] sortData_30; // @[sort.scala 28:21]
  reg [31:0] _RAND_32;
  reg [8:0] sortData_31; // @[sort.scala 28:21]
  reg [31:0] _RAND_33;
  reg [8:0] tagData_0; // @[sort.scala 29:20]
  reg [31:0] _RAND_34;
  reg [8:0] tagData_1; // @[sort.scala 29:20]
  reg [31:0] _RAND_35;
  reg [8:0] tagData_2; // @[sort.scala 29:20]
  reg [31:0] _RAND_36;
  reg [8:0] tagData_3; // @[sort.scala 29:20]
  reg [31:0] _RAND_37;
  reg [8:0] tagData_4; // @[sort.scala 29:20]
  reg [31:0] _RAND_38;
  reg [8:0] tagData_5; // @[sort.scala 29:20]
  reg [31:0] _RAND_39;
  reg [8:0] tagData_6; // @[sort.scala 29:20]
  reg [31:0] _RAND_40;
  reg [8:0] tagData_7; // @[sort.scala 29:20]
  reg [31:0] _RAND_41;
  reg [8:0] tagData_8; // @[sort.scala 29:20]
  reg [31:0] _RAND_42;
  reg [8:0] tagData_9; // @[sort.scala 29:20]
  reg [31:0] _RAND_43;
  reg [8:0] tagData_10; // @[sort.scala 29:20]
  reg [31:0] _RAND_44;
  reg [8:0] tagData_11; // @[sort.scala 29:20]
  reg [31:0] _RAND_45;
  reg [8:0] tagData_12; // @[sort.scala 29:20]
  reg [31:0] _RAND_46;
  reg [8:0] tagData_13; // @[sort.scala 29:20]
  reg [31:0] _RAND_47;
  reg [8:0] tagData_14; // @[sort.scala 29:20]
  reg [31:0] _RAND_48;
  reg [8:0] tagData_15; // @[sort.scala 29:20]
  reg [31:0] _RAND_49;
  reg [8:0] tagData_16; // @[sort.scala 29:20]
  reg [31:0] _RAND_50;
  reg [8:0] tagData_17; // @[sort.scala 29:20]
  reg [31:0] _RAND_51;
  reg [8:0] tagData_18; // @[sort.scala 29:20]
  reg [31:0] _RAND_52;
  reg [8:0] tagData_19; // @[sort.scala 29:20]
  reg [31:0] _RAND_53;
  reg [8:0] tagData_20; // @[sort.scala 29:20]
  reg [31:0] _RAND_54;
  reg [8:0] tagData_21; // @[sort.scala 29:20]
  reg [31:0] _RAND_55;
  reg [8:0] tagData_22; // @[sort.scala 29:20]
  reg [31:0] _RAND_56;
  reg [8:0] tagData_23; // @[sort.scala 29:20]
  reg [31:0] _RAND_57;
  reg [8:0] tagData_24; // @[sort.scala 29:20]
  reg [31:0] _RAND_58;
  reg [8:0] tagData_25; // @[sort.scala 29:20]
  reg [31:0] _RAND_59;
  reg [8:0] tagData_26; // @[sort.scala 29:20]
  reg [31:0] _RAND_60;
  reg [8:0] tagData_27; // @[sort.scala 29:20]
  reg [31:0] _RAND_61;
  reg [8:0] tagData_28; // @[sort.scala 29:20]
  reg [31:0] _RAND_62;
  reg [8:0] tagData_29; // @[sort.scala 29:20]
  reg [31:0] _RAND_63;
  reg [8:0] tagData_30; // @[sort.scala 29:20]
  reg [31:0] _RAND_64;
  reg [8:0] tagData_31; // @[sort.scala 29:20]
  reg [31:0] _RAND_65;
  reg [5:0] itemNumber; // @[sort.scala 30:23]
  reg [31:0] _RAND_66;
  reg [8:0] tempSortData_0; // @[sort.scala 31:25]
  reg [31:0] _RAND_67;
  reg [8:0] tempSortData_1; // @[sort.scala 31:25]
  reg [31:0] _RAND_68;
  reg [8:0] tempSortData_2; // @[sort.scala 31:25]
  reg [31:0] _RAND_69;
  reg [8:0] tempSortData_3; // @[sort.scala 31:25]
  reg [31:0] _RAND_70;
  reg [8:0] tempSortData_4; // @[sort.scala 31:25]
  reg [31:0] _RAND_71;
  reg [8:0] tempSortData_5; // @[sort.scala 31:25]
  reg [31:0] _RAND_72;
  reg [8:0] tempSortData_6; // @[sort.scala 31:25]
  reg [31:0] _RAND_73;
  reg [8:0] tempSortData_7; // @[sort.scala 31:25]
  reg [31:0] _RAND_74;
  reg [8:0] tempSortData_8; // @[sort.scala 31:25]
  reg [31:0] _RAND_75;
  reg [8:0] tempSortData_9; // @[sort.scala 31:25]
  reg [31:0] _RAND_76;
  reg [8:0] tempSortData_10; // @[sort.scala 31:25]
  reg [31:0] _RAND_77;
  reg [8:0] tempSortData_11; // @[sort.scala 31:25]
  reg [31:0] _RAND_78;
  reg [8:0] tempSortData_12; // @[sort.scala 31:25]
  reg [31:0] _RAND_79;
  reg [8:0] tempSortData_13; // @[sort.scala 31:25]
  reg [31:0] _RAND_80;
  reg [8:0] tempSortData_14; // @[sort.scala 31:25]
  reg [31:0] _RAND_81;
  reg [8:0] tempSortData_15; // @[sort.scala 31:25]
  reg [31:0] _RAND_82;
  reg [8:0] tempSortData_16; // @[sort.scala 31:25]
  reg [31:0] _RAND_83;
  reg [8:0] tempSortData_17; // @[sort.scala 31:25]
  reg [31:0] _RAND_84;
  reg [8:0] tempSortData_18; // @[sort.scala 31:25]
  reg [31:0] _RAND_85;
  reg [8:0] tempSortData_19; // @[sort.scala 31:25]
  reg [31:0] _RAND_86;
  reg [8:0] tempSortData_20; // @[sort.scala 31:25]
  reg [31:0] _RAND_87;
  reg [8:0] tempSortData_21; // @[sort.scala 31:25]
  reg [31:0] _RAND_88;
  reg [8:0] tempSortData_22; // @[sort.scala 31:25]
  reg [31:0] _RAND_89;
  reg [8:0] tempSortData_23; // @[sort.scala 31:25]
  reg [31:0] _RAND_90;
  reg [8:0] tempSortData_24; // @[sort.scala 31:25]
  reg [31:0] _RAND_91;
  reg [8:0] tempSortData_25; // @[sort.scala 31:25]
  reg [31:0] _RAND_92;
  reg [8:0] tempSortData_26; // @[sort.scala 31:25]
  reg [31:0] _RAND_93;
  reg [8:0] tempSortData_27; // @[sort.scala 31:25]
  reg [31:0] _RAND_94;
  reg [8:0] tempSortData_28; // @[sort.scala 31:25]
  reg [31:0] _RAND_95;
  reg [8:0] tempSortData_29; // @[sort.scala 31:25]
  reg [31:0] _RAND_96;
  reg [8:0] tempSortData_30; // @[sort.scala 31:25]
  reg [31:0] _RAND_97;
  reg [8:0] tempSortData_31; // @[sort.scala 31:25]
  reg [31:0] _RAND_98;
  reg [8:0] tempTagData_0; // @[sort.scala 32:24]
  reg [31:0] _RAND_99;
  reg [8:0] tempTagData_1; // @[sort.scala 32:24]
  reg [31:0] _RAND_100;
  reg [8:0] tempTagData_2; // @[sort.scala 32:24]
  reg [31:0] _RAND_101;
  reg [8:0] tempTagData_3; // @[sort.scala 32:24]
  reg [31:0] _RAND_102;
  reg [8:0] tempTagData_4; // @[sort.scala 32:24]
  reg [31:0] _RAND_103;
  reg [8:0] tempTagData_5; // @[sort.scala 32:24]
  reg [31:0] _RAND_104;
  reg [8:0] tempTagData_6; // @[sort.scala 32:24]
  reg [31:0] _RAND_105;
  reg [8:0] tempTagData_7; // @[sort.scala 32:24]
  reg [31:0] _RAND_106;
  reg [8:0] tempTagData_8; // @[sort.scala 32:24]
  reg [31:0] _RAND_107;
  reg [8:0] tempTagData_9; // @[sort.scala 32:24]
  reg [31:0] _RAND_108;
  reg [8:0] tempTagData_10; // @[sort.scala 32:24]
  reg [31:0] _RAND_109;
  reg [8:0] tempTagData_11; // @[sort.scala 32:24]
  reg [31:0] _RAND_110;
  reg [8:0] tempTagData_12; // @[sort.scala 32:24]
  reg [31:0] _RAND_111;
  reg [8:0] tempTagData_13; // @[sort.scala 32:24]
  reg [31:0] _RAND_112;
  reg [8:0] tempTagData_14; // @[sort.scala 32:24]
  reg [31:0] _RAND_113;
  reg [8:0] tempTagData_15; // @[sort.scala 32:24]
  reg [31:0] _RAND_114;
  reg [8:0] tempTagData_16; // @[sort.scala 32:24]
  reg [31:0] _RAND_115;
  reg [8:0] tempTagData_17; // @[sort.scala 32:24]
  reg [31:0] _RAND_116;
  reg [8:0] tempTagData_18; // @[sort.scala 32:24]
  reg [31:0] _RAND_117;
  reg [8:0] tempTagData_19; // @[sort.scala 32:24]
  reg [31:0] _RAND_118;
  reg [8:0] tempTagData_20; // @[sort.scala 32:24]
  reg [31:0] _RAND_119;
  reg [8:0] tempTagData_21; // @[sort.scala 32:24]
  reg [31:0] _RAND_120;
  reg [8:0] tempTagData_22; // @[sort.scala 32:24]
  reg [31:0] _RAND_121;
  reg [8:0] tempTagData_23; // @[sort.scala 32:24]
  reg [31:0] _RAND_122;
  reg [8:0] tempTagData_24; // @[sort.scala 32:24]
  reg [31:0] _RAND_123;
  reg [8:0] tempTagData_25; // @[sort.scala 32:24]
  reg [31:0] _RAND_124;
  reg [8:0] tempTagData_26; // @[sort.scala 32:24]
  reg [31:0] _RAND_125;
  reg [8:0] tempTagData_27; // @[sort.scala 32:24]
  reg [31:0] _RAND_126;
  reg [8:0] tempTagData_28; // @[sort.scala 32:24]
  reg [31:0] _RAND_127;
  reg [8:0] tempTagData_29; // @[sort.scala 32:24]
  reg [31:0] _RAND_128;
  reg [8:0] tempTagData_30; // @[sort.scala 32:24]
  reg [31:0] _RAND_129;
  reg [8:0] tempTagData_31; // @[sort.scala 32:24]
  reg [31:0] _RAND_130;
  reg [8:0] sortedSortData_0; // @[sort.scala 33:27]
  reg [31:0] _RAND_131;
  reg [8:0] sortedSortData_1; // @[sort.scala 33:27]
  reg [31:0] _RAND_132;
  reg [8:0] sortedSortData_2; // @[sort.scala 33:27]
  reg [31:0] _RAND_133;
  reg [8:0] sortedSortData_3; // @[sort.scala 33:27]
  reg [31:0] _RAND_134;
  reg [8:0] sortedSortData_4; // @[sort.scala 33:27]
  reg [31:0] _RAND_135;
  reg [8:0] sortedSortData_5; // @[sort.scala 33:27]
  reg [31:0] _RAND_136;
  reg [8:0] sortedSortData_6; // @[sort.scala 33:27]
  reg [31:0] _RAND_137;
  reg [8:0] sortedSortData_7; // @[sort.scala 33:27]
  reg [31:0] _RAND_138;
  reg [8:0] sortedSortData_8; // @[sort.scala 33:27]
  reg [31:0] _RAND_139;
  reg [8:0] sortedSortData_9; // @[sort.scala 33:27]
  reg [31:0] _RAND_140;
  reg [8:0] sortedSortData_10; // @[sort.scala 33:27]
  reg [31:0] _RAND_141;
  reg [8:0] sortedSortData_11; // @[sort.scala 33:27]
  reg [31:0] _RAND_142;
  reg [8:0] sortedSortData_12; // @[sort.scala 33:27]
  reg [31:0] _RAND_143;
  reg [8:0] sortedSortData_13; // @[sort.scala 33:27]
  reg [31:0] _RAND_144;
  reg [8:0] sortedSortData_14; // @[sort.scala 33:27]
  reg [31:0] _RAND_145;
  reg [8:0] sortedSortData_15; // @[sort.scala 33:27]
  reg [31:0] _RAND_146;
  reg [8:0] sortedSortData_16; // @[sort.scala 33:27]
  reg [31:0] _RAND_147;
  reg [8:0] sortedSortData_17; // @[sort.scala 33:27]
  reg [31:0] _RAND_148;
  reg [8:0] sortedSortData_18; // @[sort.scala 33:27]
  reg [31:0] _RAND_149;
  reg [8:0] sortedSortData_19; // @[sort.scala 33:27]
  reg [31:0] _RAND_150;
  reg [8:0] sortedSortData_20; // @[sort.scala 33:27]
  reg [31:0] _RAND_151;
  reg [8:0] sortedSortData_21; // @[sort.scala 33:27]
  reg [31:0] _RAND_152;
  reg [8:0] sortedSortData_22; // @[sort.scala 33:27]
  reg [31:0] _RAND_153;
  reg [8:0] sortedSortData_23; // @[sort.scala 33:27]
  reg [31:0] _RAND_154;
  reg [8:0] sortedSortData_24; // @[sort.scala 33:27]
  reg [31:0] _RAND_155;
  reg [8:0] sortedSortData_25; // @[sort.scala 33:27]
  reg [31:0] _RAND_156;
  reg [8:0] sortedSortData_26; // @[sort.scala 33:27]
  reg [31:0] _RAND_157;
  reg [8:0] sortedSortData_27; // @[sort.scala 33:27]
  reg [31:0] _RAND_158;
  reg [8:0] sortedSortData_28; // @[sort.scala 33:27]
  reg [31:0] _RAND_159;
  reg [8:0] sortedSortData_29; // @[sort.scala 33:27]
  reg [31:0] _RAND_160;
  reg [8:0] sortedSortData_30; // @[sort.scala 33:27]
  reg [31:0] _RAND_161;
  reg [8:0] sortedSortData_31; // @[sort.scala 33:27]
  reg [31:0] _RAND_162;
  reg [8:0] sortedTagData_0; // @[sort.scala 34:26]
  reg [31:0] _RAND_163;
  reg [8:0] sortedTagData_1; // @[sort.scala 34:26]
  reg [31:0] _RAND_164;
  reg [8:0] sortedTagData_2; // @[sort.scala 34:26]
  reg [31:0] _RAND_165;
  reg [8:0] sortedTagData_3; // @[sort.scala 34:26]
  reg [31:0] _RAND_166;
  reg [8:0] sortedTagData_4; // @[sort.scala 34:26]
  reg [31:0] _RAND_167;
  reg [8:0] sortedTagData_5; // @[sort.scala 34:26]
  reg [31:0] _RAND_168;
  reg [8:0] sortedTagData_6; // @[sort.scala 34:26]
  reg [31:0] _RAND_169;
  reg [8:0] sortedTagData_7; // @[sort.scala 34:26]
  reg [31:0] _RAND_170;
  reg [8:0] sortedTagData_8; // @[sort.scala 34:26]
  reg [31:0] _RAND_171;
  reg [8:0] sortedTagData_9; // @[sort.scala 34:26]
  reg [31:0] _RAND_172;
  reg [8:0] sortedTagData_10; // @[sort.scala 34:26]
  reg [31:0] _RAND_173;
  reg [8:0] sortedTagData_11; // @[sort.scala 34:26]
  reg [31:0] _RAND_174;
  reg [8:0] sortedTagData_12; // @[sort.scala 34:26]
  reg [31:0] _RAND_175;
  reg [8:0] sortedTagData_13; // @[sort.scala 34:26]
  reg [31:0] _RAND_176;
  reg [8:0] sortedTagData_14; // @[sort.scala 34:26]
  reg [31:0] _RAND_177;
  reg [8:0] sortedTagData_15; // @[sort.scala 34:26]
  reg [31:0] _RAND_178;
  reg [8:0] sortedTagData_16; // @[sort.scala 34:26]
  reg [31:0] _RAND_179;
  reg [8:0] sortedTagData_17; // @[sort.scala 34:26]
  reg [31:0] _RAND_180;
  reg [8:0] sortedTagData_18; // @[sort.scala 34:26]
  reg [31:0] _RAND_181;
  reg [8:0] sortedTagData_19; // @[sort.scala 34:26]
  reg [31:0] _RAND_182;
  reg [8:0] sortedTagData_20; // @[sort.scala 34:26]
  reg [31:0] _RAND_183;
  reg [8:0] sortedTagData_21; // @[sort.scala 34:26]
  reg [31:0] _RAND_184;
  reg [8:0] sortedTagData_22; // @[sort.scala 34:26]
  reg [31:0] _RAND_185;
  reg [8:0] sortedTagData_23; // @[sort.scala 34:26]
  reg [31:0] _RAND_186;
  reg [8:0] sortedTagData_24; // @[sort.scala 34:26]
  reg [31:0] _RAND_187;
  reg [8:0] sortedTagData_25; // @[sort.scala 34:26]
  reg [31:0] _RAND_188;
  reg [8:0] sortedTagData_26; // @[sort.scala 34:26]
  reg [31:0] _RAND_189;
  reg [8:0] sortedTagData_27; // @[sort.scala 34:26]
  reg [31:0] _RAND_190;
  reg [8:0] sortedTagData_28; // @[sort.scala 34:26]
  reg [31:0] _RAND_191;
  reg [8:0] sortedTagData_29; // @[sort.scala 34:26]
  reg [31:0] _RAND_192;
  reg [8:0] sortedTagData_30; // @[sort.scala 34:26]
  reg [31:0] _RAND_193;
  reg [8:0] sortedTagData_31; // @[sort.scala 34:26]
  reg [31:0] _RAND_194;
  wire  _T = ~state; // @[Conditional.scala 37:30]
  wire  _GEN_130 = io_start | state; // @[sort.scala 38:22]
  wire [5:0] _T_3 = iteration + 6'h1; // @[sort.scala 54:30]
  wire [7:0] _T_4 = itemNumber * 6'h2; // @[sort.scala 55:36]
  wire [7:0] _T_6 = _T_4 - 8'h1; // @[sort.scala 55:42]
  wire [7:0] _GEN_649 = {{2'd0}, iteration}; // @[sort.scala 55:22]
  wire  _T_7 = _GEN_649 >= _T_6; // @[sort.scala 55:22]
  wire  _T_8 = iteration < itemNumber; // @[sort.scala 58:22]
  wire  _T_11 = tempSortData_0 < sortedSortData_0; // @[sort.scala 66:34]
  wire  _T_12 = tempSortData_1 < sortedSortData_1; // @[sort.scala 66:34]
  wire  _T_13 = tempSortData_2 < sortedSortData_2; // @[sort.scala 66:34]
  wire  _T_14 = tempSortData_3 < sortedSortData_3; // @[sort.scala 66:34]
  wire  _T_15 = tempSortData_4 < sortedSortData_4; // @[sort.scala 66:34]
  wire  _T_16 = tempSortData_5 < sortedSortData_5; // @[sort.scala 66:34]
  wire  _T_17 = tempSortData_6 < sortedSortData_6; // @[sort.scala 66:34]
  wire  _T_18 = tempSortData_7 < sortedSortData_7; // @[sort.scala 66:34]
  wire  _T_19 = tempSortData_8 < sortedSortData_8; // @[sort.scala 66:34]
  wire  _T_20 = tempSortData_9 < sortedSortData_9; // @[sort.scala 66:34]
  wire  _T_21 = tempSortData_10 < sortedSortData_10; // @[sort.scala 66:34]
  wire  _T_22 = tempSortData_11 < sortedSortData_11; // @[sort.scala 66:34]
  wire  _T_23 = tempSortData_12 < sortedSortData_12; // @[sort.scala 66:34]
  wire  _T_24 = tempSortData_13 < sortedSortData_13; // @[sort.scala 66:34]
  wire  _T_25 = tempSortData_14 < sortedSortData_14; // @[sort.scala 66:34]
  wire  _T_26 = tempSortData_15 < sortedSortData_15; // @[sort.scala 66:34]
  wire  _T_27 = tempSortData_16 < sortedSortData_16; // @[sort.scala 66:34]
  wire  _T_28 = tempSortData_17 < sortedSortData_17; // @[sort.scala 66:34]
  wire  _T_29 = tempSortData_18 < sortedSortData_18; // @[sort.scala 66:34]
  wire  _T_30 = tempSortData_19 < sortedSortData_19; // @[sort.scala 66:34]
  wire  _T_31 = tempSortData_20 < sortedSortData_20; // @[sort.scala 66:34]
  wire  _T_32 = tempSortData_21 < sortedSortData_21; // @[sort.scala 66:34]
  wire  _T_33 = tempSortData_22 < sortedSortData_22; // @[sort.scala 66:34]
  wire  _T_34 = tempSortData_23 < sortedSortData_23; // @[sort.scala 66:34]
  wire  _T_35 = tempSortData_24 < sortedSortData_24; // @[sort.scala 66:34]
  wire  _T_36 = tempSortData_25 < sortedSortData_25; // @[sort.scala 66:34]
  wire  _T_37 = tempSortData_26 < sortedSortData_26; // @[sort.scala 66:34]
  wire  _T_38 = tempSortData_27 < sortedSortData_27; // @[sort.scala 66:34]
  wire  _T_39 = tempSortData_28 < sortedSortData_28; // @[sort.scala 66:34]
  wire  _T_40 = tempSortData_29 < sortedSortData_29; // @[sort.scala 66:34]
  wire  _T_41 = tempSortData_30 < sortedSortData_30; // @[sort.scala 66:34]
  wire  _T_42 = tempSortData_31 < sortedSortData_31; // @[sort.scala 66:34]
  assign io_outputs_outputData_0 = sortedSortData_0[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_1 = sortedSortData_1[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_2 = sortedSortData_2[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_3 = sortedSortData_3[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_4 = sortedSortData_4[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_5 = sortedSortData_5[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_6 = sortedSortData_6[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_7 = sortedSortData_7[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_8 = sortedSortData_8[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_9 = sortedSortData_9[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_10 = sortedSortData_10[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_11 = sortedSortData_11[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_12 = sortedSortData_12[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_13 = sortedSortData_13[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_14 = sortedSortData_14[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_15 = sortedSortData_15[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_16 = sortedSortData_16[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_17 = sortedSortData_17[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_18 = sortedSortData_18[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_19 = sortedSortData_19[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_20 = sortedSortData_20[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_21 = sortedSortData_21[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_22 = sortedSortData_22[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_23 = sortedSortData_23[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_24 = sortedSortData_24[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_25 = sortedSortData_25[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_26 = sortedSortData_26[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_27 = sortedSortData_27[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_28 = sortedSortData_28[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_29 = sortedSortData_29[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_30 = sortedSortData_30[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputData_31 = sortedSortData_31[7:0]; // @[sort.scala 83:27]
  assign io_outputs_outputTags_0 = sortedTagData_0; // @[sort.scala 84:27]
  assign io_outputs_outputTags_1 = sortedTagData_1; // @[sort.scala 84:27]
  assign io_outputs_outputTags_2 = sortedTagData_2; // @[sort.scala 84:27]
  assign io_outputs_outputTags_3 = sortedTagData_3; // @[sort.scala 84:27]
  assign io_outputs_outputTags_4 = sortedTagData_4; // @[sort.scala 84:27]
  assign io_outputs_outputTags_5 = sortedTagData_5; // @[sort.scala 84:27]
  assign io_outputs_outputTags_6 = sortedTagData_6; // @[sort.scala 84:27]
  assign io_outputs_outputTags_7 = sortedTagData_7; // @[sort.scala 84:27]
  assign io_outputs_outputTags_8 = sortedTagData_8; // @[sort.scala 84:27]
  assign io_outputs_outputTags_9 = sortedTagData_9; // @[sort.scala 84:27]
  assign io_outputs_outputTags_10 = sortedTagData_10; // @[sort.scala 84:27]
  assign io_outputs_outputTags_11 = sortedTagData_11; // @[sort.scala 84:27]
  assign io_outputs_outputTags_12 = sortedTagData_12; // @[sort.scala 84:27]
  assign io_outputs_outputTags_13 = sortedTagData_13; // @[sort.scala 84:27]
  assign io_outputs_outputTags_14 = sortedTagData_14; // @[sort.scala 84:27]
  assign io_outputs_outputTags_15 = sortedTagData_15; // @[sort.scala 84:27]
  assign io_outputs_outputTags_16 = sortedTagData_16; // @[sort.scala 84:27]
  assign io_outputs_outputTags_17 = sortedTagData_17; // @[sort.scala 84:27]
  assign io_outputs_outputTags_18 = sortedTagData_18; // @[sort.scala 84:27]
  assign io_outputs_outputTags_19 = sortedTagData_19; // @[sort.scala 84:27]
  assign io_outputs_outputTags_20 = sortedTagData_20; // @[sort.scala 84:27]
  assign io_outputs_outputTags_21 = sortedTagData_21; // @[sort.scala 84:27]
  assign io_outputs_outputTags_22 = sortedTagData_22; // @[sort.scala 84:27]
  assign io_outputs_outputTags_23 = sortedTagData_23; // @[sort.scala 84:27]
  assign io_outputs_outputTags_24 = sortedTagData_24; // @[sort.scala 84:27]
  assign io_outputs_outputTags_25 = sortedTagData_25; // @[sort.scala 84:27]
  assign io_outputs_outputTags_26 = sortedTagData_26; // @[sort.scala 84:27]
  assign io_outputs_outputTags_27 = sortedTagData_27; // @[sort.scala 84:27]
  assign io_outputs_outputTags_28 = sortedTagData_28; // @[sort.scala 84:27]
  assign io_outputs_outputTags_29 = sortedTagData_29; // @[sort.scala 84:27]
  assign io_outputs_outputTags_30 = sortedTagData_30; // @[sort.scala 84:27]
  assign io_outputs_outputTags_31 = sortedTagData_31; // @[sort.scala 84:27]
  assign io_outputs_itemNumber = itemNumber; // @[sort.scala 91:25]
  assign io_finished = ~state; // @[sort.scala 92:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  iteration = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  sortData_0 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  sortData_1 = _RAND_3[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  sortData_2 = _RAND_4[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sortData_3 = _RAND_5[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sortData_4 = _RAND_6[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sortData_5 = _RAND_7[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sortData_6 = _RAND_8[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  sortData_7 = _RAND_9[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  sortData_8 = _RAND_10[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  sortData_9 = _RAND_11[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  sortData_10 = _RAND_12[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  sortData_11 = _RAND_13[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  sortData_12 = _RAND_14[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  sortData_13 = _RAND_15[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  sortData_14 = _RAND_16[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  sortData_15 = _RAND_17[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  sortData_16 = _RAND_18[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  sortData_17 = _RAND_19[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  sortData_18 = _RAND_20[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  sortData_19 = _RAND_21[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  sortData_20 = _RAND_22[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  sortData_21 = _RAND_23[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  sortData_22 = _RAND_24[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  sortData_23 = _RAND_25[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  sortData_24 = _RAND_26[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  sortData_25 = _RAND_27[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  sortData_26 = _RAND_28[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  sortData_27 = _RAND_29[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  sortData_28 = _RAND_30[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  sortData_29 = _RAND_31[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  sortData_30 = _RAND_32[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  sortData_31 = _RAND_33[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  tagData_0 = _RAND_34[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  tagData_1 = _RAND_35[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  tagData_2 = _RAND_36[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  tagData_3 = _RAND_37[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  tagData_4 = _RAND_38[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  tagData_5 = _RAND_39[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  tagData_6 = _RAND_40[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  tagData_7 = _RAND_41[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  tagData_8 = _RAND_42[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  tagData_9 = _RAND_43[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  tagData_10 = _RAND_44[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  tagData_11 = _RAND_45[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  tagData_12 = _RAND_46[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  tagData_13 = _RAND_47[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  tagData_14 = _RAND_48[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  tagData_15 = _RAND_49[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  tagData_16 = _RAND_50[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  tagData_17 = _RAND_51[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  tagData_18 = _RAND_52[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  tagData_19 = _RAND_53[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  tagData_20 = _RAND_54[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  tagData_21 = _RAND_55[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  tagData_22 = _RAND_56[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  tagData_23 = _RAND_57[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  tagData_24 = _RAND_58[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  tagData_25 = _RAND_59[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  tagData_26 = _RAND_60[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  tagData_27 = _RAND_61[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  tagData_28 = _RAND_62[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  tagData_29 = _RAND_63[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  tagData_30 = _RAND_64[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  tagData_31 = _RAND_65[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  itemNumber = _RAND_66[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  tempSortData_0 = _RAND_67[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  tempSortData_1 = _RAND_68[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  tempSortData_2 = _RAND_69[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  tempSortData_3 = _RAND_70[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  tempSortData_4 = _RAND_71[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  tempSortData_5 = _RAND_72[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  tempSortData_6 = _RAND_73[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  tempSortData_7 = _RAND_74[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  tempSortData_8 = _RAND_75[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  tempSortData_9 = _RAND_76[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  tempSortData_10 = _RAND_77[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  tempSortData_11 = _RAND_78[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  tempSortData_12 = _RAND_79[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  tempSortData_13 = _RAND_80[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  tempSortData_14 = _RAND_81[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  tempSortData_15 = _RAND_82[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  tempSortData_16 = _RAND_83[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  tempSortData_17 = _RAND_84[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  tempSortData_18 = _RAND_85[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  tempSortData_19 = _RAND_86[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  tempSortData_20 = _RAND_87[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  tempSortData_21 = _RAND_88[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  tempSortData_22 = _RAND_89[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  tempSortData_23 = _RAND_90[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  tempSortData_24 = _RAND_91[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  tempSortData_25 = _RAND_92[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  tempSortData_26 = _RAND_93[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  tempSortData_27 = _RAND_94[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  tempSortData_28 = _RAND_95[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  tempSortData_29 = _RAND_96[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  tempSortData_30 = _RAND_97[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  tempSortData_31 = _RAND_98[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  tempTagData_0 = _RAND_99[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  tempTagData_1 = _RAND_100[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  tempTagData_2 = _RAND_101[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  tempTagData_3 = _RAND_102[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  tempTagData_4 = _RAND_103[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  tempTagData_5 = _RAND_104[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  tempTagData_6 = _RAND_105[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  tempTagData_7 = _RAND_106[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  tempTagData_8 = _RAND_107[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  tempTagData_9 = _RAND_108[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  tempTagData_10 = _RAND_109[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  tempTagData_11 = _RAND_110[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  tempTagData_12 = _RAND_111[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  tempTagData_13 = _RAND_112[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  tempTagData_14 = _RAND_113[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  tempTagData_15 = _RAND_114[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  tempTagData_16 = _RAND_115[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  tempTagData_17 = _RAND_116[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  tempTagData_18 = _RAND_117[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  tempTagData_19 = _RAND_118[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  tempTagData_20 = _RAND_119[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  tempTagData_21 = _RAND_120[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  tempTagData_22 = _RAND_121[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  tempTagData_23 = _RAND_122[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  tempTagData_24 = _RAND_123[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  tempTagData_25 = _RAND_124[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  tempTagData_26 = _RAND_125[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  tempTagData_27 = _RAND_126[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  tempTagData_28 = _RAND_127[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  tempTagData_29 = _RAND_128[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  tempTagData_30 = _RAND_129[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  tempTagData_31 = _RAND_130[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  sortedSortData_0 = _RAND_131[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  sortedSortData_1 = _RAND_132[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  sortedSortData_2 = _RAND_133[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  sortedSortData_3 = _RAND_134[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  sortedSortData_4 = _RAND_135[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  sortedSortData_5 = _RAND_136[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  sortedSortData_6 = _RAND_137[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  sortedSortData_7 = _RAND_138[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  sortedSortData_8 = _RAND_139[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  sortedSortData_9 = _RAND_140[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  sortedSortData_10 = _RAND_141[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  sortedSortData_11 = _RAND_142[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  sortedSortData_12 = _RAND_143[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  sortedSortData_13 = _RAND_144[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  sortedSortData_14 = _RAND_145[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  sortedSortData_15 = _RAND_146[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  sortedSortData_16 = _RAND_147[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  sortedSortData_17 = _RAND_148[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  sortedSortData_18 = _RAND_149[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  sortedSortData_19 = _RAND_150[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  sortedSortData_20 = _RAND_151[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  sortedSortData_21 = _RAND_152[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  sortedSortData_22 = _RAND_153[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  sortedSortData_23 = _RAND_154[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  sortedSortData_24 = _RAND_155[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  sortedSortData_25 = _RAND_156[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  sortedSortData_26 = _RAND_157[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  sortedSortData_27 = _RAND_158[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  sortedSortData_28 = _RAND_159[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  sortedSortData_29 = _RAND_160[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  sortedSortData_30 = _RAND_161[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  sortedSortData_31 = _RAND_162[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  sortedTagData_0 = _RAND_163[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  sortedTagData_1 = _RAND_164[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  sortedTagData_2 = _RAND_165[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  sortedTagData_3 = _RAND_166[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  sortedTagData_4 = _RAND_167[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  sortedTagData_5 = _RAND_168[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  sortedTagData_6 = _RAND_169[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  sortedTagData_7 = _RAND_170[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  sortedTagData_8 = _RAND_171[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  sortedTagData_9 = _RAND_172[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  sortedTagData_10 = _RAND_173[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  sortedTagData_11 = _RAND_174[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  sortedTagData_12 = _RAND_175[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  sortedTagData_13 = _RAND_176[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  sortedTagData_14 = _RAND_177[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  sortedTagData_15 = _RAND_178[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  sortedTagData_16 = _RAND_179[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  sortedTagData_17 = _RAND_180[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  sortedTagData_18 = _RAND_181[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  sortedTagData_19 = _RAND_182[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  sortedTagData_20 = _RAND_183[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  sortedTagData_21 = _RAND_184[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  sortedTagData_22 = _RAND_185[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  sortedTagData_23 = _RAND_186[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  sortedTagData_24 = _RAND_187[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  sortedTagData_25 = _RAND_188[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  sortedTagData_26 = _RAND_189[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  sortedTagData_27 = _RAND_190[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  sortedTagData_28 = _RAND_191[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  sortedTagData_29 = _RAND_192[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  sortedTagData_30 = _RAND_193[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  sortedTagData_31 = _RAND_194[8:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else if (_T) begin
      state <= _GEN_130;
    end else if (state) begin
      if (_T_7) begin
        state <= 1'h0;
      end
    end
    if (_T) begin
      if (io_start) begin
        iteration <= 6'h0;
      end
    end else if (state) begin
      iteration <= _T_3;
    end
    if (_T) begin
      if (io_start) begin
        sortData_0 <= {{3'd0}, io_inputs_depths_0};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_1 <= {{3'd0}, io_inputs_depths_1};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_2 <= {{3'd0}, io_inputs_depths_2};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_3 <= {{3'd0}, io_inputs_depths_3};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_4 <= {{3'd0}, io_inputs_depths_4};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_5 <= {{3'd0}, io_inputs_depths_5};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_6 <= {{3'd0}, io_inputs_depths_6};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_7 <= {{3'd0}, io_inputs_depths_7};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_8 <= {{3'd0}, io_inputs_depths_8};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_9 <= {{3'd0}, io_inputs_depths_9};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_10 <= {{3'd0}, io_inputs_depths_10};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_11 <= {{3'd0}, io_inputs_depths_11};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_12 <= {{3'd0}, io_inputs_depths_12};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_13 <= {{3'd0}, io_inputs_depths_13};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_14 <= {{3'd0}, io_inputs_depths_14};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_15 <= {{3'd0}, io_inputs_depths_15};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_16 <= {{3'd0}, io_inputs_depths_16};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_17 <= {{3'd0}, io_inputs_depths_17};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_18 <= {{3'd0}, io_inputs_depths_18};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_19 <= {{3'd0}, io_inputs_depths_19};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_20 <= {{3'd0}, io_inputs_depths_20};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_21 <= {{3'd0}, io_inputs_depths_21};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_22 <= {{3'd0}, io_inputs_depths_22};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_23 <= {{3'd0}, io_inputs_depths_23};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_24 <= {{3'd0}, io_inputs_depths_24};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_25 <= {{3'd0}, io_inputs_depths_25};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_26 <= {{3'd0}, io_inputs_depths_26};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_27 <= {{3'd0}, io_inputs_depths_27};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_28 <= {{3'd0}, io_inputs_depths_28};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_29 <= {{3'd0}, io_inputs_depths_29};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_30 <= {{3'd0}, io_inputs_depths_30};
      end
    end
    if (_T) begin
      if (io_start) begin
        sortData_31 <= {{3'd0}, io_inputs_depths_31};
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_0 <= io_inputs_characters_0;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_1 <= io_inputs_characters_1;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_2 <= io_inputs_characters_2;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_3 <= io_inputs_characters_3;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_4 <= io_inputs_characters_4;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_5 <= io_inputs_characters_5;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_6 <= io_inputs_characters_6;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_7 <= io_inputs_characters_7;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_8 <= io_inputs_characters_8;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_9 <= io_inputs_characters_9;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_10 <= io_inputs_characters_10;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_11 <= io_inputs_characters_11;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_12 <= io_inputs_characters_12;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_13 <= io_inputs_characters_13;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_14 <= io_inputs_characters_14;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_15 <= io_inputs_characters_15;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_16 <= io_inputs_characters_16;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_17 <= io_inputs_characters_17;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_18 <= io_inputs_characters_18;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_19 <= io_inputs_characters_19;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_20 <= io_inputs_characters_20;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_21 <= io_inputs_characters_21;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_22 <= io_inputs_characters_22;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_23 <= io_inputs_characters_23;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_24 <= io_inputs_characters_24;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_25 <= io_inputs_characters_25;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_26 <= io_inputs_characters_26;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_27 <= io_inputs_characters_27;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_28 <= io_inputs_characters_28;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_29 <= io_inputs_characters_29;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_30 <= io_inputs_characters_30;
      end
    end
    if (_T) begin
      if (io_start) begin
        tagData_31 <= io_inputs_characters_31;
      end
    end
    if (_T) begin
      if (io_start) begin
        itemNumber <= io_inputs_validCharacters;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_0 <= 9'h100;
      end
    end else if (state) begin
      if (_T_8) begin
        if (5'h1f == iteration[4:0]) begin
          tempSortData_0 <= sortData_31;
        end else if (5'h1e == iteration[4:0]) begin
          tempSortData_0 <= sortData_30;
        end else if (5'h1d == iteration[4:0]) begin
          tempSortData_0 <= sortData_29;
        end else if (5'h1c == iteration[4:0]) begin
          tempSortData_0 <= sortData_28;
        end else if (5'h1b == iteration[4:0]) begin
          tempSortData_0 <= sortData_27;
        end else if (5'h1a == iteration[4:0]) begin
          tempSortData_0 <= sortData_26;
        end else if (5'h19 == iteration[4:0]) begin
          tempSortData_0 <= sortData_25;
        end else if (5'h18 == iteration[4:0]) begin
          tempSortData_0 <= sortData_24;
        end else if (5'h17 == iteration[4:0]) begin
          tempSortData_0 <= sortData_23;
        end else if (5'h16 == iteration[4:0]) begin
          tempSortData_0 <= sortData_22;
        end else if (5'h15 == iteration[4:0]) begin
          tempSortData_0 <= sortData_21;
        end else if (5'h14 == iteration[4:0]) begin
          tempSortData_0 <= sortData_20;
        end else if (5'h13 == iteration[4:0]) begin
          tempSortData_0 <= sortData_19;
        end else if (5'h12 == iteration[4:0]) begin
          tempSortData_0 <= sortData_18;
        end else if (5'h11 == iteration[4:0]) begin
          tempSortData_0 <= sortData_17;
        end else if (5'h10 == iteration[4:0]) begin
          tempSortData_0 <= sortData_16;
        end else if (5'hf == iteration[4:0]) begin
          tempSortData_0 <= sortData_15;
        end else if (5'he == iteration[4:0]) begin
          tempSortData_0 <= sortData_14;
        end else if (5'hd == iteration[4:0]) begin
          tempSortData_0 <= sortData_13;
        end else if (5'hc == iteration[4:0]) begin
          tempSortData_0 <= sortData_12;
        end else if (5'hb == iteration[4:0]) begin
          tempSortData_0 <= sortData_11;
        end else if (5'ha == iteration[4:0]) begin
          tempSortData_0 <= sortData_10;
        end else if (5'h9 == iteration[4:0]) begin
          tempSortData_0 <= sortData_9;
        end else if (5'h8 == iteration[4:0]) begin
          tempSortData_0 <= sortData_8;
        end else if (5'h7 == iteration[4:0]) begin
          tempSortData_0 <= sortData_7;
        end else if (5'h6 == iteration[4:0]) begin
          tempSortData_0 <= sortData_6;
        end else if (5'h5 == iteration[4:0]) begin
          tempSortData_0 <= sortData_5;
        end else if (5'h4 == iteration[4:0]) begin
          tempSortData_0 <= sortData_4;
        end else if (5'h3 == iteration[4:0]) begin
          tempSortData_0 <= sortData_3;
        end else if (5'h2 == iteration[4:0]) begin
          tempSortData_0 <= sortData_2;
        end else if (5'h1 == iteration[4:0]) begin
          tempSortData_0 <= sortData_1;
        end else begin
          tempSortData_0 <= sortData_0;
        end
      end else begin
        tempSortData_0 <= 9'h100;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_1 <= 9'h100;
      end
    end else if (state) begin
      if (_T_11) begin
        tempSortData_1 <= sortedSortData_0;
      end else begin
        tempSortData_1 <= tempSortData_0;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_2 <= 9'h100;
      end
    end else if (state) begin
      if (_T_12) begin
        tempSortData_2 <= sortedSortData_1;
      end else begin
        tempSortData_2 <= tempSortData_1;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_3 <= 9'h100;
      end
    end else if (state) begin
      if (_T_13) begin
        tempSortData_3 <= sortedSortData_2;
      end else begin
        tempSortData_3 <= tempSortData_2;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_4 <= 9'h100;
      end
    end else if (state) begin
      if (_T_14) begin
        tempSortData_4 <= sortedSortData_3;
      end else begin
        tempSortData_4 <= tempSortData_3;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_5 <= 9'h100;
      end
    end else if (state) begin
      if (_T_15) begin
        tempSortData_5 <= sortedSortData_4;
      end else begin
        tempSortData_5 <= tempSortData_4;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_6 <= 9'h100;
      end
    end else if (state) begin
      if (_T_16) begin
        tempSortData_6 <= sortedSortData_5;
      end else begin
        tempSortData_6 <= tempSortData_5;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_7 <= 9'h100;
      end
    end else if (state) begin
      if (_T_17) begin
        tempSortData_7 <= sortedSortData_6;
      end else begin
        tempSortData_7 <= tempSortData_6;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_8 <= 9'h100;
      end
    end else if (state) begin
      if (_T_18) begin
        tempSortData_8 <= sortedSortData_7;
      end else begin
        tempSortData_8 <= tempSortData_7;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_9 <= 9'h100;
      end
    end else if (state) begin
      if (_T_19) begin
        tempSortData_9 <= sortedSortData_8;
      end else begin
        tempSortData_9 <= tempSortData_8;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_10 <= 9'h100;
      end
    end else if (state) begin
      if (_T_20) begin
        tempSortData_10 <= sortedSortData_9;
      end else begin
        tempSortData_10 <= tempSortData_9;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_11 <= 9'h100;
      end
    end else if (state) begin
      if (_T_21) begin
        tempSortData_11 <= sortedSortData_10;
      end else begin
        tempSortData_11 <= tempSortData_10;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_12 <= 9'h100;
      end
    end else if (state) begin
      if (_T_22) begin
        tempSortData_12 <= sortedSortData_11;
      end else begin
        tempSortData_12 <= tempSortData_11;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_13 <= 9'h100;
      end
    end else if (state) begin
      if (_T_23) begin
        tempSortData_13 <= sortedSortData_12;
      end else begin
        tempSortData_13 <= tempSortData_12;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_14 <= 9'h100;
      end
    end else if (state) begin
      if (_T_24) begin
        tempSortData_14 <= sortedSortData_13;
      end else begin
        tempSortData_14 <= tempSortData_13;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_15 <= 9'h100;
      end
    end else if (state) begin
      if (_T_25) begin
        tempSortData_15 <= sortedSortData_14;
      end else begin
        tempSortData_15 <= tempSortData_14;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_16 <= 9'h100;
      end
    end else if (state) begin
      if (_T_26) begin
        tempSortData_16 <= sortedSortData_15;
      end else begin
        tempSortData_16 <= tempSortData_15;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_17 <= 9'h100;
      end
    end else if (state) begin
      if (_T_27) begin
        tempSortData_17 <= sortedSortData_16;
      end else begin
        tempSortData_17 <= tempSortData_16;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_18 <= 9'h100;
      end
    end else if (state) begin
      if (_T_28) begin
        tempSortData_18 <= sortedSortData_17;
      end else begin
        tempSortData_18 <= tempSortData_17;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_19 <= 9'h100;
      end
    end else if (state) begin
      if (_T_29) begin
        tempSortData_19 <= sortedSortData_18;
      end else begin
        tempSortData_19 <= tempSortData_18;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_20 <= 9'h100;
      end
    end else if (state) begin
      if (_T_30) begin
        tempSortData_20 <= sortedSortData_19;
      end else begin
        tempSortData_20 <= tempSortData_19;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_21 <= 9'h100;
      end
    end else if (state) begin
      if (_T_31) begin
        tempSortData_21 <= sortedSortData_20;
      end else begin
        tempSortData_21 <= tempSortData_20;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_22 <= 9'h100;
      end
    end else if (state) begin
      if (_T_32) begin
        tempSortData_22 <= sortedSortData_21;
      end else begin
        tempSortData_22 <= tempSortData_21;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_23 <= 9'h100;
      end
    end else if (state) begin
      if (_T_33) begin
        tempSortData_23 <= sortedSortData_22;
      end else begin
        tempSortData_23 <= tempSortData_22;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_24 <= 9'h100;
      end
    end else if (state) begin
      if (_T_34) begin
        tempSortData_24 <= sortedSortData_23;
      end else begin
        tempSortData_24 <= tempSortData_23;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_25 <= 9'h100;
      end
    end else if (state) begin
      if (_T_35) begin
        tempSortData_25 <= sortedSortData_24;
      end else begin
        tempSortData_25 <= tempSortData_24;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_26 <= 9'h100;
      end
    end else if (state) begin
      if (_T_36) begin
        tempSortData_26 <= sortedSortData_25;
      end else begin
        tempSortData_26 <= tempSortData_25;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_27 <= 9'h100;
      end
    end else if (state) begin
      if (_T_37) begin
        tempSortData_27 <= sortedSortData_26;
      end else begin
        tempSortData_27 <= tempSortData_26;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_28 <= 9'h100;
      end
    end else if (state) begin
      if (_T_38) begin
        tempSortData_28 <= sortedSortData_27;
      end else begin
        tempSortData_28 <= tempSortData_27;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_29 <= 9'h100;
      end
    end else if (state) begin
      if (_T_39) begin
        tempSortData_29 <= sortedSortData_28;
      end else begin
        tempSortData_29 <= tempSortData_28;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_30 <= 9'h100;
      end
    end else if (state) begin
      if (_T_40) begin
        tempSortData_30 <= sortedSortData_29;
      end else begin
        tempSortData_30 <= tempSortData_29;
      end
    end
    if (_T) begin
      if (io_start) begin
        tempSortData_31 <= 9'h100;
      end
    end else if (state) begin
      if (_T_41) begin
        tempSortData_31 <= sortedSortData_30;
      end else begin
        tempSortData_31 <= tempSortData_30;
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_8) begin
          if (5'h1f == iteration[4:0]) begin
            tempTagData_0 <= tagData_31;
          end else if (5'h1e == iteration[4:0]) begin
            tempTagData_0 <= tagData_30;
          end else if (5'h1d == iteration[4:0]) begin
            tempTagData_0 <= tagData_29;
          end else if (5'h1c == iteration[4:0]) begin
            tempTagData_0 <= tagData_28;
          end else if (5'h1b == iteration[4:0]) begin
            tempTagData_0 <= tagData_27;
          end else if (5'h1a == iteration[4:0]) begin
            tempTagData_0 <= tagData_26;
          end else if (5'h19 == iteration[4:0]) begin
            tempTagData_0 <= tagData_25;
          end else if (5'h18 == iteration[4:0]) begin
            tempTagData_0 <= tagData_24;
          end else if (5'h17 == iteration[4:0]) begin
            tempTagData_0 <= tagData_23;
          end else if (5'h16 == iteration[4:0]) begin
            tempTagData_0 <= tagData_22;
          end else if (5'h15 == iteration[4:0]) begin
            tempTagData_0 <= tagData_21;
          end else if (5'h14 == iteration[4:0]) begin
            tempTagData_0 <= tagData_20;
          end else if (5'h13 == iteration[4:0]) begin
            tempTagData_0 <= tagData_19;
          end else if (5'h12 == iteration[4:0]) begin
            tempTagData_0 <= tagData_18;
          end else if (5'h11 == iteration[4:0]) begin
            tempTagData_0 <= tagData_17;
          end else if (5'h10 == iteration[4:0]) begin
            tempTagData_0 <= tagData_16;
          end else if (5'hf == iteration[4:0]) begin
            tempTagData_0 <= tagData_15;
          end else if (5'he == iteration[4:0]) begin
            tempTagData_0 <= tagData_14;
          end else if (5'hd == iteration[4:0]) begin
            tempTagData_0 <= tagData_13;
          end else if (5'hc == iteration[4:0]) begin
            tempTagData_0 <= tagData_12;
          end else if (5'hb == iteration[4:0]) begin
            tempTagData_0 <= tagData_11;
          end else if (5'ha == iteration[4:0]) begin
            tempTagData_0 <= tagData_10;
          end else if (5'h9 == iteration[4:0]) begin
            tempTagData_0 <= tagData_9;
          end else if (5'h8 == iteration[4:0]) begin
            tempTagData_0 <= tagData_8;
          end else if (5'h7 == iteration[4:0]) begin
            tempTagData_0 <= tagData_7;
          end else if (5'h6 == iteration[4:0]) begin
            tempTagData_0 <= tagData_6;
          end else if (5'h5 == iteration[4:0]) begin
            tempTagData_0 <= tagData_5;
          end else if (5'h4 == iteration[4:0]) begin
            tempTagData_0 <= tagData_4;
          end else if (5'h3 == iteration[4:0]) begin
            tempTagData_0 <= tagData_3;
          end else if (5'h2 == iteration[4:0]) begin
            tempTagData_0 <= tagData_2;
          end else if (5'h1 == iteration[4:0]) begin
            tempTagData_0 <= tagData_1;
          end else begin
            tempTagData_0 <= tagData_0;
          end
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_11) begin
          tempTagData_1 <= sortedTagData_0;
        end else begin
          tempTagData_1 <= tempTagData_0;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_12) begin
          tempTagData_2 <= sortedTagData_1;
        end else begin
          tempTagData_2 <= tempTagData_1;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_13) begin
          tempTagData_3 <= sortedTagData_2;
        end else begin
          tempTagData_3 <= tempTagData_2;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_14) begin
          tempTagData_4 <= sortedTagData_3;
        end else begin
          tempTagData_4 <= tempTagData_3;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_15) begin
          tempTagData_5 <= sortedTagData_4;
        end else begin
          tempTagData_5 <= tempTagData_4;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_16) begin
          tempTagData_6 <= sortedTagData_5;
        end else begin
          tempTagData_6 <= tempTagData_5;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_17) begin
          tempTagData_7 <= sortedTagData_6;
        end else begin
          tempTagData_7 <= tempTagData_6;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_18) begin
          tempTagData_8 <= sortedTagData_7;
        end else begin
          tempTagData_8 <= tempTagData_7;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_19) begin
          tempTagData_9 <= sortedTagData_8;
        end else begin
          tempTagData_9 <= tempTagData_8;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_20) begin
          tempTagData_10 <= sortedTagData_9;
        end else begin
          tempTagData_10 <= tempTagData_9;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_21) begin
          tempTagData_11 <= sortedTagData_10;
        end else begin
          tempTagData_11 <= tempTagData_10;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_22) begin
          tempTagData_12 <= sortedTagData_11;
        end else begin
          tempTagData_12 <= tempTagData_11;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_23) begin
          tempTagData_13 <= sortedTagData_12;
        end else begin
          tempTagData_13 <= tempTagData_12;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_24) begin
          tempTagData_14 <= sortedTagData_13;
        end else begin
          tempTagData_14 <= tempTagData_13;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_25) begin
          tempTagData_15 <= sortedTagData_14;
        end else begin
          tempTagData_15 <= tempTagData_14;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_26) begin
          tempTagData_16 <= sortedTagData_15;
        end else begin
          tempTagData_16 <= tempTagData_15;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_27) begin
          tempTagData_17 <= sortedTagData_16;
        end else begin
          tempTagData_17 <= tempTagData_16;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_28) begin
          tempTagData_18 <= sortedTagData_17;
        end else begin
          tempTagData_18 <= tempTagData_17;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_29) begin
          tempTagData_19 <= sortedTagData_18;
        end else begin
          tempTagData_19 <= tempTagData_18;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_30) begin
          tempTagData_20 <= sortedTagData_19;
        end else begin
          tempTagData_20 <= tempTagData_19;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_31) begin
          tempTagData_21 <= sortedTagData_20;
        end else begin
          tempTagData_21 <= tempTagData_20;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_32) begin
          tempTagData_22 <= sortedTagData_21;
        end else begin
          tempTagData_22 <= tempTagData_21;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_33) begin
          tempTagData_23 <= sortedTagData_22;
        end else begin
          tempTagData_23 <= tempTagData_22;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_34) begin
          tempTagData_24 <= sortedTagData_23;
        end else begin
          tempTagData_24 <= tempTagData_23;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_35) begin
          tempTagData_25 <= sortedTagData_24;
        end else begin
          tempTagData_25 <= tempTagData_24;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_36) begin
          tempTagData_26 <= sortedTagData_25;
        end else begin
          tempTagData_26 <= tempTagData_25;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_37) begin
          tempTagData_27 <= sortedTagData_26;
        end else begin
          tempTagData_27 <= tempTagData_26;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_38) begin
          tempTagData_28 <= sortedTagData_27;
        end else begin
          tempTagData_28 <= tempTagData_27;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_39) begin
          tempTagData_29 <= sortedTagData_28;
        end else begin
          tempTagData_29 <= tempTagData_28;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_40) begin
          tempTagData_30 <= sortedTagData_29;
        end else begin
          tempTagData_30 <= tempTagData_29;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_41) begin
          tempTagData_31 <= sortedTagData_30;
        end else begin
          tempTagData_31 <= tempTagData_30;
        end
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_0 <= 9'h100;
      end
    end else if (state) begin
      if (_T_11) begin
        sortedSortData_0 <= tempSortData_0;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_1 <= 9'h100;
      end
    end else if (state) begin
      if (_T_12) begin
        sortedSortData_1 <= tempSortData_1;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_2 <= 9'h100;
      end
    end else if (state) begin
      if (_T_13) begin
        sortedSortData_2 <= tempSortData_2;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_3 <= 9'h100;
      end
    end else if (state) begin
      if (_T_14) begin
        sortedSortData_3 <= tempSortData_3;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_4 <= 9'h100;
      end
    end else if (state) begin
      if (_T_15) begin
        sortedSortData_4 <= tempSortData_4;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_5 <= 9'h100;
      end
    end else if (state) begin
      if (_T_16) begin
        sortedSortData_5 <= tempSortData_5;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_6 <= 9'h100;
      end
    end else if (state) begin
      if (_T_17) begin
        sortedSortData_6 <= tempSortData_6;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_7 <= 9'h100;
      end
    end else if (state) begin
      if (_T_18) begin
        sortedSortData_7 <= tempSortData_7;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_8 <= 9'h100;
      end
    end else if (state) begin
      if (_T_19) begin
        sortedSortData_8 <= tempSortData_8;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_9 <= 9'h100;
      end
    end else if (state) begin
      if (_T_20) begin
        sortedSortData_9 <= tempSortData_9;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_10 <= 9'h100;
      end
    end else if (state) begin
      if (_T_21) begin
        sortedSortData_10 <= tempSortData_10;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_11 <= 9'h100;
      end
    end else if (state) begin
      if (_T_22) begin
        sortedSortData_11 <= tempSortData_11;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_12 <= 9'h100;
      end
    end else if (state) begin
      if (_T_23) begin
        sortedSortData_12 <= tempSortData_12;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_13 <= 9'h100;
      end
    end else if (state) begin
      if (_T_24) begin
        sortedSortData_13 <= tempSortData_13;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_14 <= 9'h100;
      end
    end else if (state) begin
      if (_T_25) begin
        sortedSortData_14 <= tempSortData_14;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_15 <= 9'h100;
      end
    end else if (state) begin
      if (_T_26) begin
        sortedSortData_15 <= tempSortData_15;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_16 <= 9'h100;
      end
    end else if (state) begin
      if (_T_27) begin
        sortedSortData_16 <= tempSortData_16;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_17 <= 9'h100;
      end
    end else if (state) begin
      if (_T_28) begin
        sortedSortData_17 <= tempSortData_17;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_18 <= 9'h100;
      end
    end else if (state) begin
      if (_T_29) begin
        sortedSortData_18 <= tempSortData_18;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_19 <= 9'h100;
      end
    end else if (state) begin
      if (_T_30) begin
        sortedSortData_19 <= tempSortData_19;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_20 <= 9'h100;
      end
    end else if (state) begin
      if (_T_31) begin
        sortedSortData_20 <= tempSortData_20;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_21 <= 9'h100;
      end
    end else if (state) begin
      if (_T_32) begin
        sortedSortData_21 <= tempSortData_21;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_22 <= 9'h100;
      end
    end else if (state) begin
      if (_T_33) begin
        sortedSortData_22 <= tempSortData_22;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_23 <= 9'h100;
      end
    end else if (state) begin
      if (_T_34) begin
        sortedSortData_23 <= tempSortData_23;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_24 <= 9'h100;
      end
    end else if (state) begin
      if (_T_35) begin
        sortedSortData_24 <= tempSortData_24;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_25 <= 9'h100;
      end
    end else if (state) begin
      if (_T_36) begin
        sortedSortData_25 <= tempSortData_25;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_26 <= 9'h100;
      end
    end else if (state) begin
      if (_T_37) begin
        sortedSortData_26 <= tempSortData_26;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_27 <= 9'h100;
      end
    end else if (state) begin
      if (_T_38) begin
        sortedSortData_27 <= tempSortData_27;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_28 <= 9'h100;
      end
    end else if (state) begin
      if (_T_39) begin
        sortedSortData_28 <= tempSortData_28;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_29 <= 9'h100;
      end
    end else if (state) begin
      if (_T_40) begin
        sortedSortData_29 <= tempSortData_29;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_30 <= 9'h100;
      end
    end else if (state) begin
      if (_T_41) begin
        sortedSortData_30 <= tempSortData_30;
      end
    end
    if (_T) begin
      if (io_start) begin
        sortedSortData_31 <= 9'h100;
      end
    end else if (state) begin
      if (_T_42) begin
        sortedSortData_31 <= tempSortData_31;
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_11) begin
          sortedTagData_0 <= tempTagData_0;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_12) begin
          sortedTagData_1 <= tempTagData_1;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_13) begin
          sortedTagData_2 <= tempTagData_2;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_14) begin
          sortedTagData_3 <= tempTagData_3;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_15) begin
          sortedTagData_4 <= tempTagData_4;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_16) begin
          sortedTagData_5 <= tempTagData_5;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_17) begin
          sortedTagData_6 <= tempTagData_6;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_18) begin
          sortedTagData_7 <= tempTagData_7;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_19) begin
          sortedTagData_8 <= tempTagData_8;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_20) begin
          sortedTagData_9 <= tempTagData_9;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_21) begin
          sortedTagData_10 <= tempTagData_10;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_22) begin
          sortedTagData_11 <= tempTagData_11;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_23) begin
          sortedTagData_12 <= tempTagData_12;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_24) begin
          sortedTagData_13 <= tempTagData_13;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_25) begin
          sortedTagData_14 <= tempTagData_14;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_26) begin
          sortedTagData_15 <= tempTagData_15;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_27) begin
          sortedTagData_16 <= tempTagData_16;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_28) begin
          sortedTagData_17 <= tempTagData_17;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_29) begin
          sortedTagData_18 <= tempTagData_18;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_30) begin
          sortedTagData_19 <= tempTagData_19;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_31) begin
          sortedTagData_20 <= tempTagData_20;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_32) begin
          sortedTagData_21 <= tempTagData_21;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_33) begin
          sortedTagData_22 <= tempTagData_22;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_34) begin
          sortedTagData_23 <= tempTagData_23;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_35) begin
          sortedTagData_24 <= tempTagData_24;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_36) begin
          sortedTagData_25 <= tempTagData_25;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_37) begin
          sortedTagData_26 <= tempTagData_26;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_38) begin
          sortedTagData_27 <= tempTagData_27;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_39) begin
          sortedTagData_28 <= tempTagData_28;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_40) begin
          sortedTagData_29 <= tempTagData_29;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_41) begin
          sortedTagData_30 <= tempTagData_30;
        end
      end
    end
    if (!(_T)) begin
      if (state) begin
        if (_T_42) begin
          sortedTagData_31 <= tempTagData_31;
        end
      end
    end
  end
endmodule
module treeNormalizer(
  input        clock,
  input        reset,
  input        io_start,
  input  [7:0] io_inputs_outputData_0,
  input  [7:0] io_inputs_outputData_1,
  input  [7:0] io_inputs_outputData_2,
  input  [7:0] io_inputs_outputData_3,
  input  [7:0] io_inputs_outputData_4,
  input  [7:0] io_inputs_outputData_5,
  input  [7:0] io_inputs_outputData_6,
  input  [7:0] io_inputs_outputData_7,
  input  [7:0] io_inputs_outputData_8,
  input  [7:0] io_inputs_outputData_9,
  input  [7:0] io_inputs_outputData_10,
  input  [7:0] io_inputs_outputData_11,
  input  [7:0] io_inputs_outputData_12,
  input  [7:0] io_inputs_outputData_13,
  input  [7:0] io_inputs_outputData_14,
  input  [7:0] io_inputs_outputData_15,
  input  [7:0] io_inputs_outputData_16,
  input  [7:0] io_inputs_outputData_17,
  input  [7:0] io_inputs_outputData_18,
  input  [7:0] io_inputs_outputData_19,
  input  [7:0] io_inputs_outputData_20,
  input  [7:0] io_inputs_outputData_21,
  input  [7:0] io_inputs_outputData_22,
  input  [7:0] io_inputs_outputData_23,
  input  [7:0] io_inputs_outputData_24,
  input  [7:0] io_inputs_outputData_25,
  input  [7:0] io_inputs_outputData_26,
  input  [7:0] io_inputs_outputData_27,
  input  [7:0] io_inputs_outputData_28,
  input  [7:0] io_inputs_outputData_29,
  input  [7:0] io_inputs_outputData_30,
  input  [7:0] io_inputs_outputData_31,
  input  [8:0] io_inputs_outputTags_0,
  input  [8:0] io_inputs_outputTags_1,
  input  [8:0] io_inputs_outputTags_2,
  input  [8:0] io_inputs_outputTags_3,
  input  [8:0] io_inputs_outputTags_4,
  input  [8:0] io_inputs_outputTags_5,
  input  [8:0] io_inputs_outputTags_6,
  input  [8:0] io_inputs_outputTags_7,
  input  [8:0] io_inputs_outputTags_8,
  input  [8:0] io_inputs_outputTags_9,
  input  [8:0] io_inputs_outputTags_10,
  input  [8:0] io_inputs_outputTags_11,
  input  [8:0] io_inputs_outputTags_12,
  input  [8:0] io_inputs_outputTags_13,
  input  [8:0] io_inputs_outputTags_14,
  input  [8:0] io_inputs_outputTags_15,
  input  [8:0] io_inputs_outputTags_16,
  input  [8:0] io_inputs_outputTags_17,
  input  [8:0] io_inputs_outputTags_18,
  input  [8:0] io_inputs_outputTags_19,
  input  [8:0] io_inputs_outputTags_20,
  input  [8:0] io_inputs_outputTags_21,
  input  [8:0] io_inputs_outputTags_22,
  input  [8:0] io_inputs_outputTags_23,
  input  [8:0] io_inputs_outputTags_24,
  input  [8:0] io_inputs_outputTags_25,
  input  [8:0] io_inputs_outputTags_26,
  input  [8:0] io_inputs_outputTags_27,
  input  [8:0] io_inputs_outputTags_28,
  input  [8:0] io_inputs_outputTags_29,
  input  [8:0] io_inputs_outputTags_30,
  input  [8:0] io_inputs_outputTags_31,
  input  [5:0] io_inputs_itemNumber,
  output [8:0] io_outputs_charactersOut_0,
  output [8:0] io_outputs_charactersOut_1,
  output [8:0] io_outputs_charactersOut_2,
  output [8:0] io_outputs_charactersOut_3,
  output [8:0] io_outputs_charactersOut_4,
  output [8:0] io_outputs_charactersOut_5,
  output [8:0] io_outputs_charactersOut_6,
  output [8:0] io_outputs_charactersOut_7,
  output [8:0] io_outputs_charactersOut_8,
  output [8:0] io_outputs_charactersOut_9,
  output [8:0] io_outputs_charactersOut_10,
  output [8:0] io_outputs_charactersOut_11,
  output [8:0] io_outputs_charactersOut_12,
  output [8:0] io_outputs_charactersOut_13,
  output [8:0] io_outputs_charactersOut_14,
  output [8:0] io_outputs_charactersOut_15,
  output [8:0] io_outputs_charactersOut_16,
  output [8:0] io_outputs_charactersOut_17,
  output [8:0] io_outputs_charactersOut_18,
  output [8:0] io_outputs_charactersOut_19,
  output [8:0] io_outputs_charactersOut_20,
  output [8:0] io_outputs_charactersOut_21,
  output [8:0] io_outputs_charactersOut_22,
  output [8:0] io_outputs_charactersOut_23,
  output [8:0] io_outputs_charactersOut_24,
  output [8:0] io_outputs_charactersOut_25,
  output [8:0] io_outputs_charactersOut_26,
  output [8:0] io_outputs_charactersOut_27,
  output [8:0] io_outputs_charactersOut_28,
  output [8:0] io_outputs_charactersOut_29,
  output [8:0] io_outputs_charactersOut_30,
  output [8:0] io_outputs_charactersOut_31,
  output [7:0] io_outputs_depthsOut_0,
  output [7:0] io_outputs_depthsOut_1,
  output [7:0] io_outputs_depthsOut_2,
  output [7:0] io_outputs_depthsOut_3,
  output [7:0] io_outputs_depthsOut_4,
  output [7:0] io_outputs_depthsOut_5,
  output [7:0] io_outputs_depthsOut_6,
  output [7:0] io_outputs_depthsOut_7,
  output [7:0] io_outputs_depthsOut_8,
  output [7:0] io_outputs_depthsOut_9,
  output [7:0] io_outputs_depthsOut_10,
  output [7:0] io_outputs_depthsOut_11,
  output [7:0] io_outputs_depthsOut_12,
  output [7:0] io_outputs_depthsOut_13,
  output [7:0] io_outputs_depthsOut_14,
  output [7:0] io_outputs_depthsOut_15,
  output [7:0] io_outputs_depthsOut_16,
  output [7:0] io_outputs_depthsOut_17,
  output [7:0] io_outputs_depthsOut_18,
  output [7:0] io_outputs_depthsOut_19,
  output [7:0] io_outputs_depthsOut_20,
  output [7:0] io_outputs_depthsOut_21,
  output [7:0] io_outputs_depthsOut_22,
  output [7:0] io_outputs_depthsOut_23,
  output [7:0] io_outputs_depthsOut_24,
  output [7:0] io_outputs_depthsOut_25,
  output [7:0] io_outputs_depthsOut_26,
  output [7:0] io_outputs_depthsOut_27,
  output [7:0] io_outputs_depthsOut_28,
  output [7:0] io_outputs_depthsOut_29,
  output [7:0] io_outputs_depthsOut_30,
  output [7:0] io_outputs_depthsOut_31,
  output [8:0] io_outputs_validNodesOut,
  output       io_finished
);
  reg [1:0] state; // @[treeNormalizer.scala 37:22]
  reg [31:0] _RAND_0;
  reg [7:0] depthsOut_0; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_1;
  reg [7:0] depthsOut_1; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_2;
  reg [7:0] depthsOut_2; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_3;
  reg [7:0] depthsOut_3; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_4;
  reg [7:0] depthsOut_4; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_5;
  reg [7:0] depthsOut_5; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_6;
  reg [7:0] depthsOut_6; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_7;
  reg [7:0] depthsOut_7; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_8;
  reg [7:0] depthsOut_8; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_9;
  reg [7:0] depthsOut_9; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_10;
  reg [7:0] depthsOut_10; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_11;
  reg [7:0] depthsOut_11; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_12;
  reg [7:0] depthsOut_12; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_13;
  reg [7:0] depthsOut_13; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_14;
  reg [7:0] depthsOut_14; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_15;
  reg [7:0] depthsOut_15; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_16;
  reg [7:0] depthsOut_16; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_17;
  reg [7:0] depthsOut_17; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_18;
  reg [7:0] depthsOut_18; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_19;
  reg [7:0] depthsOut_19; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_20;
  reg [7:0] depthsOut_20; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_21;
  reg [7:0] depthsOut_21; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_22;
  reg [7:0] depthsOut_22; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_23;
  reg [7:0] depthsOut_23; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_24;
  reg [7:0] depthsOut_24; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_25;
  reg [7:0] depthsOut_25; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_26;
  reg [7:0] depthsOut_26; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_27;
  reg [7:0] depthsOut_27; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_28;
  reg [7:0] depthsOut_28; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_29;
  reg [7:0] depthsOut_29; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_30;
  reg [7:0] depthsOut_30; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_31;
  reg [7:0] depthsOut_31; // @[treeNormalizer.scala 39:22]
  reg [31:0] _RAND_32;
  reg [5:0] charactersAtDepth_0; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_33;
  reg [5:0] charactersAtDepth_1; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_34;
  reg [5:0] charactersAtDepth_2; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_35;
  reg [5:0] charactersAtDepth_3; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_36;
  reg [5:0] charactersAtDepth_4; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_37;
  reg [5:0] charactersAtDepth_5; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_38;
  reg [5:0] charactersAtDepth_6; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_39;
  reg [5:0] charactersAtDepth_7; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_40;
  reg [5:0] charactersAtDepth_8; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_41;
  reg [5:0] charactersAtDepth_9; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_42;
  reg [5:0] charactersAtDepth_10; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_43;
  reg [5:0] charactersAtDepth_11; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_44;
  reg [5:0] charactersAtDepth_12; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_45;
  reg [5:0] charactersAtDepth_13; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_46;
  reg [5:0] charactersAtDepth_14; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_47;
  reg [5:0] charactersAtDepth_15; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_48;
  reg [5:0] charactersAtDepth_16; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_49;
  reg [5:0] charactersAtDepth_17; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_50;
  reg [5:0] charactersAtDepth_18; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_51;
  reg [5:0] charactersAtDepth_19; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_52;
  reg [5:0] charactersAtDepth_20; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_53;
  reg [5:0] charactersAtDepth_21; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_54;
  reg [5:0] charactersAtDepth_22; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_55;
  reg [5:0] charactersAtDepth_23; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_56;
  reg [5:0] charactersAtDepth_24; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_57;
  reg [5:0] charactersAtDepth_25; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_58;
  reg [5:0] charactersAtDepth_26; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_59;
  reg [5:0] charactersAtDepth_27; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_60;
  reg [5:0] charactersAtDepth_28; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_61;
  reg [5:0] charactersAtDepth_29; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_62;
  reg [5:0] charactersAtDepth_30; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_63;
  reg [5:0] charactersAtDepth_31; // @[treeNormalizer.scala 65:30]
  reg [31:0] _RAND_64;
  wire [36:0] _T_1 = {$signed(charactersAtDepth_0), 31'h0}; // @[treeNormalizer.scala 80:49]
  wire [32:0] subtractCharacters_0 = _T_1[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 80:25]
  wire [32:0] _GEN_653 = {{27{charactersAtDepth_1[5]}},charactersAtDepth_1}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_4 = $signed(subtractCharacters_0) + $signed(_GEN_653); // @[treeNormalizer.scala 82:64]
  wire [62:0] _T_5 = {$signed(_T_4), 30'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_1 = _T_5[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_655 = {{27{charactersAtDepth_2[5]}},charactersAtDepth_2}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_8 = $signed(subtractCharacters_1) + $signed(_GEN_655); // @[treeNormalizer.scala 82:64]
  wire [61:0] _T_9 = {$signed(_T_8), 29'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_2 = _T_9[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_657 = {{27{charactersAtDepth_3[5]}},charactersAtDepth_3}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_12 = $signed(subtractCharacters_2) + $signed(_GEN_657); // @[treeNormalizer.scala 82:64]
  wire [60:0] _T_13 = {$signed(_T_12), 28'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_3 = _T_13[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_659 = {{27{charactersAtDepth_4[5]}},charactersAtDepth_4}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_16 = $signed(subtractCharacters_3) + $signed(_GEN_659); // @[treeNormalizer.scala 82:64]
  wire [59:0] _T_17 = {$signed(_T_16), 27'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_4 = _T_17[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_661 = {{27{charactersAtDepth_5[5]}},charactersAtDepth_5}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_20 = $signed(subtractCharacters_4) + $signed(_GEN_661); // @[treeNormalizer.scala 82:64]
  wire [58:0] _T_21 = {$signed(_T_20), 26'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_5 = _T_21[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_663 = {{27{charactersAtDepth_6[5]}},charactersAtDepth_6}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_24 = $signed(subtractCharacters_5) + $signed(_GEN_663); // @[treeNormalizer.scala 82:64]
  wire [57:0] _T_25 = {$signed(_T_24), 25'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_6 = _T_25[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_665 = {{27{charactersAtDepth_7[5]}},charactersAtDepth_7}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_28 = $signed(subtractCharacters_6) + $signed(_GEN_665); // @[treeNormalizer.scala 82:64]
  wire [56:0] _T_29 = {$signed(_T_28), 24'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_7 = _T_29[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_667 = {{27{charactersAtDepth_8[5]}},charactersAtDepth_8}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_32 = $signed(subtractCharacters_7) + $signed(_GEN_667); // @[treeNormalizer.scala 82:64]
  wire [55:0] _T_33 = {$signed(_T_32), 23'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_8 = _T_33[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_669 = {{27{charactersAtDepth_9[5]}},charactersAtDepth_9}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_36 = $signed(subtractCharacters_8) + $signed(_GEN_669); // @[treeNormalizer.scala 82:64]
  wire [54:0] _T_37 = {$signed(_T_36), 22'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_9 = _T_37[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_671 = {{27{charactersAtDepth_10[5]}},charactersAtDepth_10}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_40 = $signed(subtractCharacters_9) + $signed(_GEN_671); // @[treeNormalizer.scala 82:64]
  wire [53:0] _T_41 = {$signed(_T_40), 21'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_10 = _T_41[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_673 = {{27{charactersAtDepth_11[5]}},charactersAtDepth_11}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_44 = $signed(subtractCharacters_10) + $signed(_GEN_673); // @[treeNormalizer.scala 82:64]
  wire [52:0] _T_45 = {$signed(_T_44), 20'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_11 = _T_45[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_675 = {{27{charactersAtDepth_12[5]}},charactersAtDepth_12}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_48 = $signed(subtractCharacters_11) + $signed(_GEN_675); // @[treeNormalizer.scala 82:64]
  wire [51:0] _T_49 = {$signed(_T_48), 19'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_12 = _T_49[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_677 = {{27{charactersAtDepth_13[5]}},charactersAtDepth_13}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_52 = $signed(subtractCharacters_12) + $signed(_GEN_677); // @[treeNormalizer.scala 82:64]
  wire [50:0] _T_53 = {$signed(_T_52), 18'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_13 = _T_53[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_679 = {{27{charactersAtDepth_14[5]}},charactersAtDepth_14}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_56 = $signed(subtractCharacters_13) + $signed(_GEN_679); // @[treeNormalizer.scala 82:64]
  wire [49:0] _T_57 = {$signed(_T_56), 17'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_14 = _T_57[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_681 = {{27{charactersAtDepth_15[5]}},charactersAtDepth_15}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_60 = $signed(subtractCharacters_14) + $signed(_GEN_681); // @[treeNormalizer.scala 82:64]
  wire [48:0] _T_61 = {$signed(_T_60), 16'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_15 = _T_61[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_683 = {{27{charactersAtDepth_16[5]}},charactersAtDepth_16}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_64 = $signed(subtractCharacters_15) + $signed(_GEN_683); // @[treeNormalizer.scala 82:64]
  wire [47:0] _T_65 = {$signed(_T_64), 15'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_16 = _T_65[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_685 = {{27{charactersAtDepth_17[5]}},charactersAtDepth_17}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_68 = $signed(subtractCharacters_16) + $signed(_GEN_685); // @[treeNormalizer.scala 82:64]
  wire [46:0] _T_69 = {$signed(_T_68), 14'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_17 = _T_69[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_687 = {{27{charactersAtDepth_18[5]}},charactersAtDepth_18}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_72 = $signed(subtractCharacters_17) + $signed(_GEN_687); // @[treeNormalizer.scala 82:64]
  wire [45:0] _T_73 = {$signed(_T_72), 13'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_18 = _T_73[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_689 = {{27{charactersAtDepth_19[5]}},charactersAtDepth_19}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_76 = $signed(subtractCharacters_18) + $signed(_GEN_689); // @[treeNormalizer.scala 82:64]
  wire [44:0] _T_77 = {$signed(_T_76), 12'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_19 = _T_77[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_691 = {{27{charactersAtDepth_20[5]}},charactersAtDepth_20}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_80 = $signed(subtractCharacters_19) + $signed(_GEN_691); // @[treeNormalizer.scala 82:64]
  wire [43:0] _T_81 = {$signed(_T_80), 11'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_20 = _T_81[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_693 = {{27{charactersAtDepth_21[5]}},charactersAtDepth_21}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_84 = $signed(subtractCharacters_20) + $signed(_GEN_693); // @[treeNormalizer.scala 82:64]
  wire [42:0] _T_85 = {$signed(_T_84), 10'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_21 = _T_85[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_695 = {{27{charactersAtDepth_22[5]}},charactersAtDepth_22}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_88 = $signed(subtractCharacters_21) + $signed(_GEN_695); // @[treeNormalizer.scala 82:64]
  wire [41:0] _T_89 = {$signed(_T_88), 9'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_22 = _T_89[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_697 = {{27{charactersAtDepth_23[5]}},charactersAtDepth_23}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_92 = $signed(subtractCharacters_22) + $signed(_GEN_697); // @[treeNormalizer.scala 82:64]
  wire [40:0] _T_93 = {$signed(_T_92), 8'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_23 = _T_93[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_699 = {{27{charactersAtDepth_24[5]}},charactersAtDepth_24}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_96 = $signed(subtractCharacters_23) + $signed(_GEN_699); // @[treeNormalizer.scala 82:64]
  wire [39:0] _T_97 = {$signed(_T_96), 7'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_24 = _T_97[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_701 = {{27{charactersAtDepth_25[5]}},charactersAtDepth_25}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_100 = $signed(subtractCharacters_24) + $signed(_GEN_701); // @[treeNormalizer.scala 82:64]
  wire [38:0] _T_101 = {$signed(_T_100), 6'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_25 = _T_101[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_703 = {{27{charactersAtDepth_26[5]}},charactersAtDepth_26}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_104 = $signed(subtractCharacters_25) + $signed(_GEN_703); // @[treeNormalizer.scala 82:64]
  wire [37:0] _T_105 = {$signed(_T_104), 5'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_26 = _T_105[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_705 = {{27{charactersAtDepth_27[5]}},charactersAtDepth_27}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_108 = $signed(subtractCharacters_26) + $signed(_GEN_705); // @[treeNormalizer.scala 82:64]
  wire [36:0] _T_109 = {$signed(_T_108), 4'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_27 = _T_109[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_707 = {{27{charactersAtDepth_28[5]}},charactersAtDepth_28}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_112 = $signed(subtractCharacters_27) + $signed(_GEN_707); // @[treeNormalizer.scala 82:64]
  wire [35:0] _T_113 = {$signed(_T_112), 3'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_28 = _T_113[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_709 = {{27{charactersAtDepth_29[5]}},charactersAtDepth_29}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_116 = $signed(subtractCharacters_28) + $signed(_GEN_709); // @[treeNormalizer.scala 82:64]
  wire [34:0] _T_117 = {$signed(_T_116), 2'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_29 = _T_117[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_711 = {{27{charactersAtDepth_30[5]}},charactersAtDepth_30}; // @[treeNormalizer.scala 82:64]
  wire [32:0] _T_120 = $signed(subtractCharacters_29) + $signed(_GEN_711); // @[treeNormalizer.scala 82:64]
  wire [33:0] _T_121 = {$signed(_T_120), 1'h0}; // @[treeNormalizer.scala 84:7]
  wire [32:0] subtractCharacters_30 = _T_121[32:0]; // @[treeNormalizer.scala 71:32 treeNormalizer.scala 82:31]
  wire [32:0] _GEN_713 = {{27{charactersAtDepth_31[5]}},charactersAtDepth_31}; // @[treeNormalizer.scala 82:64]
  wire [32:0] subtractCharacters_31 = $signed(subtractCharacters_30) + $signed(_GEN_713); // @[treeNormalizer.scala 82:64]
  wire [33:0] _GEN_714 = {{1{subtractCharacters_31[32]}},subtractCharacters_31}; // @[treeNormalizer.scala 86:43]
  wire [33:0] _T_129 = 34'sh100000000 - $signed(_GEN_714); // @[treeNormalizer.scala 86:43]
  reg [5:0] iteration; // @[treeNormalizer.scala 90:22]
  reg [31:0] _RAND_65;
  wire  _T_130 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_132 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_36 = 5'h1 == iteration[4:0] ? io_inputs_outputData_1 : io_inputs_outputData_0; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_37 = 5'h2 == iteration[4:0] ? io_inputs_outputData_2 : _GEN_36; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_38 = 5'h3 == iteration[4:0] ? io_inputs_outputData_3 : _GEN_37; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_39 = 5'h4 == iteration[4:0] ? io_inputs_outputData_4 : _GEN_38; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_40 = 5'h5 == iteration[4:0] ? io_inputs_outputData_5 : _GEN_39; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_41 = 5'h6 == iteration[4:0] ? io_inputs_outputData_6 : _GEN_40; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_42 = 5'h7 == iteration[4:0] ? io_inputs_outputData_7 : _GEN_41; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_43 = 5'h8 == iteration[4:0] ? io_inputs_outputData_8 : _GEN_42; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_44 = 5'h9 == iteration[4:0] ? io_inputs_outputData_9 : _GEN_43; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_45 = 5'ha == iteration[4:0] ? io_inputs_outputData_10 : _GEN_44; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_46 = 5'hb == iteration[4:0] ? io_inputs_outputData_11 : _GEN_45; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_47 = 5'hc == iteration[4:0] ? io_inputs_outputData_12 : _GEN_46; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_48 = 5'hd == iteration[4:0] ? io_inputs_outputData_13 : _GEN_47; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_49 = 5'he == iteration[4:0] ? io_inputs_outputData_14 : _GEN_48; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_50 = 5'hf == iteration[4:0] ? io_inputs_outputData_15 : _GEN_49; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_51 = 5'h10 == iteration[4:0] ? io_inputs_outputData_16 : _GEN_50; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_52 = 5'h11 == iteration[4:0] ? io_inputs_outputData_17 : _GEN_51; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_53 = 5'h12 == iteration[4:0] ? io_inputs_outputData_18 : _GEN_52; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_54 = 5'h13 == iteration[4:0] ? io_inputs_outputData_19 : _GEN_53; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_55 = 5'h14 == iteration[4:0] ? io_inputs_outputData_20 : _GEN_54; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_56 = 5'h15 == iteration[4:0] ? io_inputs_outputData_21 : _GEN_55; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_57 = 5'h16 == iteration[4:0] ? io_inputs_outputData_22 : _GEN_56; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_58 = 5'h17 == iteration[4:0] ? io_inputs_outputData_23 : _GEN_57; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_59 = 5'h18 == iteration[4:0] ? io_inputs_outputData_24 : _GEN_58; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_60 = 5'h19 == iteration[4:0] ? io_inputs_outputData_25 : _GEN_59; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_61 = 5'h1a == iteration[4:0] ? io_inputs_outputData_26 : _GEN_60; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_62 = 5'h1b == iteration[4:0] ? io_inputs_outputData_27 : _GEN_61; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_63 = 5'h1c == iteration[4:0] ? io_inputs_outputData_28 : _GEN_62; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_64 = 5'h1d == iteration[4:0] ? io_inputs_outputData_29 : _GEN_63; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_65 = 5'h1e == iteration[4:0] ? io_inputs_outputData_30 : _GEN_64; // @[treeNormalizer.scala 108:32]
  wire [7:0] _GEN_66 = 5'h1f == iteration[4:0] ? io_inputs_outputData_31 : _GEN_65; // @[treeNormalizer.scala 108:32]
  wire  _T_134 = _GEN_66 > 8'h20; // @[treeNormalizer.scala 108:32]
  wire [5:0] _T_137 = $signed(charactersAtDepth_31) + 6'sh1; // @[treeNormalizer.scala 111:11]
  wire [5:0] _GEN_68 = 5'h1 == iteration[4:0] ? $signed(charactersAtDepth_1) : $signed(charactersAtDepth_0); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_69 = 5'h2 == iteration[4:0] ? $signed(charactersAtDepth_2) : $signed(_GEN_68); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_70 = 5'h3 == iteration[4:0] ? $signed(charactersAtDepth_3) : $signed(_GEN_69); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_71 = 5'h4 == iteration[4:0] ? $signed(charactersAtDepth_4) : $signed(_GEN_70); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_72 = 5'h5 == iteration[4:0] ? $signed(charactersAtDepth_5) : $signed(_GEN_71); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_73 = 5'h6 == iteration[4:0] ? $signed(charactersAtDepth_6) : $signed(_GEN_72); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_74 = 5'h7 == iteration[4:0] ? $signed(charactersAtDepth_7) : $signed(_GEN_73); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_75 = 5'h8 == iteration[4:0] ? $signed(charactersAtDepth_8) : $signed(_GEN_74); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_76 = 5'h9 == iteration[4:0] ? $signed(charactersAtDepth_9) : $signed(_GEN_75); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_77 = 5'ha == iteration[4:0] ? $signed(charactersAtDepth_10) : $signed(_GEN_76); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_78 = 5'hb == iteration[4:0] ? $signed(charactersAtDepth_11) : $signed(_GEN_77); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_79 = 5'hc == iteration[4:0] ? $signed(charactersAtDepth_12) : $signed(_GEN_78); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_80 = 5'hd == iteration[4:0] ? $signed(charactersAtDepth_13) : $signed(_GEN_79); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_81 = 5'he == iteration[4:0] ? $signed(charactersAtDepth_14) : $signed(_GEN_80); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_82 = 5'hf == iteration[4:0] ? $signed(charactersAtDepth_15) : $signed(_GEN_81); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_83 = 5'h10 == iteration[4:0] ? $signed(charactersAtDepth_16) : $signed(_GEN_82); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_84 = 5'h11 == iteration[4:0] ? $signed(charactersAtDepth_17) : $signed(_GEN_83); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_85 = 5'h12 == iteration[4:0] ? $signed(charactersAtDepth_18) : $signed(_GEN_84); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_86 = 5'h13 == iteration[4:0] ? $signed(charactersAtDepth_19) : $signed(_GEN_85); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_87 = 5'h14 == iteration[4:0] ? $signed(charactersAtDepth_20) : $signed(_GEN_86); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_88 = 5'h15 == iteration[4:0] ? $signed(charactersAtDepth_21) : $signed(_GEN_87); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_89 = 5'h16 == iteration[4:0] ? $signed(charactersAtDepth_22) : $signed(_GEN_88); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_90 = 5'h17 == iteration[4:0] ? $signed(charactersAtDepth_23) : $signed(_GEN_89); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_91 = 5'h18 == iteration[4:0] ? $signed(charactersAtDepth_24) : $signed(_GEN_90); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_92 = 5'h19 == iteration[4:0] ? $signed(charactersAtDepth_25) : $signed(_GEN_91); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_93 = 5'h1a == iteration[4:0] ? $signed(charactersAtDepth_26) : $signed(_GEN_92); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_94 = 5'h1b == iteration[4:0] ? $signed(charactersAtDepth_27) : $signed(_GEN_93); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_95 = 5'h1c == iteration[4:0] ? $signed(charactersAtDepth_28) : $signed(_GEN_94); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_96 = 5'h1d == iteration[4:0] ? $signed(charactersAtDepth_29) : $signed(_GEN_95); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_97 = 5'h1e == iteration[4:0] ? $signed(charactersAtDepth_30) : $signed(_GEN_96); // @[treeNormalizer.scala 113:70]
  wire [5:0] _GEN_98 = 5'h1f == iteration[4:0] ? $signed(charactersAtDepth_31) : $signed(_GEN_97); // @[treeNormalizer.scala 113:70]
  wire [5:0] _T_142 = $signed(_GEN_98) + 6'sh1; // @[treeNormalizer.scala 113:70]
  wire [5:0] _T_144 = iteration + 6'h1; // @[treeNormalizer.scala 116:30]
  wire [8:0] validNodesIn = {{3'd0}, io_inputs_itemNumber}; // @[treeNormalizer.scala 43:9 treeNormalizer.scala 58:18]
  wire [8:0] _GEN_715 = {{3'd0}, _T_144}; // @[treeNormalizer.scala 118:26]
  wire  _T_147 = _GEN_715 >= validNodesIn; // @[treeNormalizer.scala 118:26]
  wire  _T_150 = _T_144 >= 6'h20; // @[treeNormalizer.scala 118:63]
  wire  _T_151 = _T_147 | _T_150; // @[treeNormalizer.scala 118:43]
  wire  _T_152 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire [32:0] freeCharacters = _T_129[32:0]; // @[treeNormalizer.scala 77:28 treeNormalizer.scala 79:18 treeNormalizer.scala 86:18]
  wire  _T_156 = $signed(freeCharacters) >= 33'sh0; // @[treeNormalizer.scala 128:29]
  wire [7:0] _T_162 = _GEN_66 - 8'h1; // @[treeNormalizer.scala 131:55]
  wire [5:0] _T_166 = iteration - 6'h1; // @[treeNormalizer.scala 136:30]
  wire  _T_167 = iteration == 6'h0; // @[treeNormalizer.scala 137:22]
  assign io_outputs_charactersOut_0 = io_inputs_outputTags_0; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_1 = io_inputs_outputTags_1; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_2 = io_inputs_outputTags_2; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_3 = io_inputs_outputTags_3; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_4 = io_inputs_outputTags_4; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_5 = io_inputs_outputTags_5; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_6 = io_inputs_outputTags_6; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_7 = io_inputs_outputTags_7; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_8 = io_inputs_outputTags_8; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_9 = io_inputs_outputTags_9; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_10 = io_inputs_outputTags_10; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_11 = io_inputs_outputTags_11; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_12 = io_inputs_outputTags_12; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_13 = io_inputs_outputTags_13; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_14 = io_inputs_outputTags_14; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_15 = io_inputs_outputTags_15; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_16 = io_inputs_outputTags_16; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_17 = io_inputs_outputTags_17; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_18 = io_inputs_outputTags_18; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_19 = io_inputs_outputTags_19; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_20 = io_inputs_outputTags_20; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_21 = io_inputs_outputTags_21; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_22 = io_inputs_outputTags_22; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_23 = io_inputs_outputTags_23; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_24 = io_inputs_outputTags_24; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_25 = io_inputs_outputTags_25; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_26 = io_inputs_outputTags_26; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_27 = io_inputs_outputTags_27; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_28 = io_inputs_outputTags_28; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_29 = io_inputs_outputTags_29; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_30 = io_inputs_outputTags_30; // @[treeNormalizer.scala 143:28]
  assign io_outputs_charactersOut_31 = io_inputs_outputTags_31; // @[treeNormalizer.scala 143:28]
  assign io_outputs_depthsOut_0 = depthsOut_0; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_1 = depthsOut_1; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_2 = depthsOut_2; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_3 = depthsOut_3; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_4 = depthsOut_4; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_5 = depthsOut_5; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_6 = depthsOut_6; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_7 = depthsOut_7; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_8 = depthsOut_8; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_9 = depthsOut_9; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_10 = depthsOut_10; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_11 = depthsOut_11; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_12 = depthsOut_12; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_13 = depthsOut_13; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_14 = depthsOut_14; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_15 = depthsOut_15; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_16 = depthsOut_16; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_17 = depthsOut_17; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_18 = depthsOut_18; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_19 = depthsOut_19; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_20 = depthsOut_20; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_21 = depthsOut_21; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_22 = depthsOut_22; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_23 = depthsOut_23; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_24 = depthsOut_24; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_25 = depthsOut_25; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_26 = depthsOut_26; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_27 = depthsOut_27; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_28 = depthsOut_28; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_29 = depthsOut_29; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_30 = depthsOut_30; // @[treeNormalizer.scala 144:24]
  assign io_outputs_depthsOut_31 = depthsOut_31; // @[treeNormalizer.scala 144:24]
  assign io_outputs_validNodesOut = {{3'd0}, io_inputs_itemNumber}; // @[treeNormalizer.scala 145:28]
  assign io_finished = state == 2'h0; // @[treeNormalizer.scala 146:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  depthsOut_0 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  depthsOut_1 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  depthsOut_2 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  depthsOut_3 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  depthsOut_4 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  depthsOut_5 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  depthsOut_6 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  depthsOut_7 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  depthsOut_8 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  depthsOut_9 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  depthsOut_10 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  depthsOut_11 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  depthsOut_12 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  depthsOut_13 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  depthsOut_14 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  depthsOut_15 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  depthsOut_16 = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  depthsOut_17 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  depthsOut_18 = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  depthsOut_19 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  depthsOut_20 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  depthsOut_21 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  depthsOut_22 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  depthsOut_23 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  depthsOut_24 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  depthsOut_25 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  depthsOut_26 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  depthsOut_27 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  depthsOut_28 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  depthsOut_29 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  depthsOut_30 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  depthsOut_31 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  charactersAtDepth_0 = _RAND_33[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  charactersAtDepth_1 = _RAND_34[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  charactersAtDepth_2 = _RAND_35[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  charactersAtDepth_3 = _RAND_36[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  charactersAtDepth_4 = _RAND_37[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  charactersAtDepth_5 = _RAND_38[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  charactersAtDepth_6 = _RAND_39[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  charactersAtDepth_7 = _RAND_40[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  charactersAtDepth_8 = _RAND_41[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  charactersAtDepth_9 = _RAND_42[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  charactersAtDepth_10 = _RAND_43[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  charactersAtDepth_11 = _RAND_44[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  charactersAtDepth_12 = _RAND_45[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  charactersAtDepth_13 = _RAND_46[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  charactersAtDepth_14 = _RAND_47[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  charactersAtDepth_15 = _RAND_48[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  charactersAtDepth_16 = _RAND_49[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  charactersAtDepth_17 = _RAND_50[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  charactersAtDepth_18 = _RAND_51[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  charactersAtDepth_19 = _RAND_52[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  charactersAtDepth_20 = _RAND_53[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  charactersAtDepth_21 = _RAND_54[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  charactersAtDepth_22 = _RAND_55[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  charactersAtDepth_23 = _RAND_56[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  charactersAtDepth_24 = _RAND_57[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  charactersAtDepth_25 = _RAND_58[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  charactersAtDepth_26 = _RAND_59[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  charactersAtDepth_27 = _RAND_60[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  charactersAtDepth_28 = _RAND_61[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  charactersAtDepth_29 = _RAND_62[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  charactersAtDepth_30 = _RAND_63[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  charactersAtDepth_31 = _RAND_64[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  iteration = _RAND_65[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T_130) begin
      if (io_start) begin
        state <= 2'h2;
      end
    end else if (_T_132) begin
      if (_T_151) begin
        state <= 2'h1;
      end
    end else if (_T_152) begin
      if (_T_167) begin
        state <= 2'h0;
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h0 == iteration[4:0]) begin
              depthsOut_0 <= 8'h20;
            end
          end else if (5'h0 == iteration[4:0]) begin
            if (5'h1f == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_31;
            end else if (5'h1e == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_30;
            end else if (5'h1d == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_29;
            end else if (5'h1c == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_28;
            end else if (5'h1b == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_27;
            end else if (5'h1a == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_26;
            end else if (5'h19 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_25;
            end else if (5'h18 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_24;
            end else if (5'h17 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_23;
            end else if (5'h16 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_22;
            end else if (5'h15 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_21;
            end else if (5'h14 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_20;
            end else if (5'h13 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_19;
            end else if (5'h12 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_18;
            end else if (5'h11 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_17;
            end else if (5'h10 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_16;
            end else if (5'hf == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_15;
            end else if (5'he == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_14;
            end else if (5'hd == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_13;
            end else if (5'hc == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_12;
            end else if (5'hb == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_11;
            end else if (5'ha == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_10;
            end else if (5'h9 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_9;
            end else if (5'h8 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_8;
            end else if (5'h7 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_7;
            end else if (5'h6 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_6;
            end else if (5'h5 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_5;
            end else if (5'h4 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_4;
            end else if (5'h3 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_3;
            end else if (5'h2 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_2;
            end else if (5'h1 == iteration[4:0]) begin
              depthsOut_0 <= io_inputs_outputData_1;
            end else begin
              depthsOut_0 <= io_inputs_outputData_0;
            end
          end else if (_T_156) begin
            if (5'h0 == iteration[4:0]) begin
              if (5'h1f == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_31;
              end else if (5'h1e == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_30;
              end else if (5'h1d == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_29;
              end else if (5'h1c == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_28;
              end else if (5'h1b == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_27;
              end else if (5'h1a == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_26;
              end else if (5'h19 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_25;
              end else if (5'h18 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_24;
              end else if (5'h17 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_23;
              end else if (5'h16 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_22;
              end else if (5'h15 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_21;
              end else if (5'h14 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_20;
              end else if (5'h13 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_19;
              end else if (5'h12 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_18;
              end else if (5'h11 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_17;
              end else if (5'h10 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_16;
              end else if (5'hf == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_15;
              end else if (5'he == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_14;
              end else if (5'hd == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_13;
              end else if (5'hc == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_12;
              end else if (5'hb == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_11;
              end else if (5'ha == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_10;
              end else if (5'h9 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_9;
              end else if (5'h8 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_8;
              end else if (5'h7 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_7;
              end else if (5'h6 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_6;
              end else if (5'h5 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_5;
              end else if (5'h4 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_4;
              end else if (5'h3 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_3;
              end else if (5'h2 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_2;
              end else if (5'h1 == iteration[4:0]) begin
                depthsOut_0 <= io_inputs_outputData_1;
              end else begin
                depthsOut_0 <= io_inputs_outputData_0;
              end
            end
          end else if (5'h0 == iteration[4:0]) begin
            depthsOut_0 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h1 == iteration[4:0]) begin
              depthsOut_1 <= 8'h20;
            end
          end else if (5'h1 == iteration[4:0]) begin
            if (5'h1f == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_31;
            end else if (5'h1e == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_30;
            end else if (5'h1d == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_29;
            end else if (5'h1c == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_28;
            end else if (5'h1b == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_27;
            end else if (5'h1a == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_26;
            end else if (5'h19 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_25;
            end else if (5'h18 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_24;
            end else if (5'h17 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_23;
            end else if (5'h16 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_22;
            end else if (5'h15 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_21;
            end else if (5'h14 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_20;
            end else if (5'h13 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_19;
            end else if (5'h12 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_18;
            end else if (5'h11 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_17;
            end else if (5'h10 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_16;
            end else if (5'hf == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_15;
            end else if (5'he == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_14;
            end else if (5'hd == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_13;
            end else if (5'hc == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_12;
            end else if (5'hb == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_11;
            end else if (5'ha == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_10;
            end else if (5'h9 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_9;
            end else if (5'h8 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_8;
            end else if (5'h7 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_7;
            end else if (5'h6 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_6;
            end else if (5'h5 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_5;
            end else if (5'h4 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_4;
            end else if (5'h3 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_3;
            end else if (5'h2 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_2;
            end else if (5'h1 == iteration[4:0]) begin
              depthsOut_1 <= io_inputs_outputData_1;
            end else begin
              depthsOut_1 <= io_inputs_outputData_0;
            end
          end else if (_T_156) begin
            if (5'h1 == iteration[4:0]) begin
              if (5'h1f == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_31;
              end else if (5'h1e == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_30;
              end else if (5'h1d == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_29;
              end else if (5'h1c == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_28;
              end else if (5'h1b == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_27;
              end else if (5'h1a == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_26;
              end else if (5'h19 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_25;
              end else if (5'h18 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_24;
              end else if (5'h17 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_23;
              end else if (5'h16 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_22;
              end else if (5'h15 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_21;
              end else if (5'h14 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_20;
              end else if (5'h13 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_19;
              end else if (5'h12 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_18;
              end else if (5'h11 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_17;
              end else if (5'h10 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_16;
              end else if (5'hf == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_15;
              end else if (5'he == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_14;
              end else if (5'hd == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_13;
              end else if (5'hc == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_12;
              end else if (5'hb == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_11;
              end else if (5'ha == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_10;
              end else if (5'h9 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_9;
              end else if (5'h8 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_8;
              end else if (5'h7 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_7;
              end else if (5'h6 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_6;
              end else if (5'h5 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_5;
              end else if (5'h4 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_4;
              end else if (5'h3 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_3;
              end else if (5'h2 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_2;
              end else if (5'h1 == iteration[4:0]) begin
                depthsOut_1 <= io_inputs_outputData_1;
              end else begin
                depthsOut_1 <= io_inputs_outputData_0;
              end
            end
          end else if (5'h1 == iteration[4:0]) begin
            depthsOut_1 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h2 == iteration[4:0]) begin
              depthsOut_2 <= 8'h20;
            end
          end else if (5'h2 == iteration[4:0]) begin
            depthsOut_2 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h2 == iteration[4:0]) begin
              depthsOut_2 <= _GEN_66;
            end
          end else if (5'h2 == iteration[4:0]) begin
            depthsOut_2 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h3 == iteration[4:0]) begin
              depthsOut_3 <= 8'h20;
            end
          end else if (5'h3 == iteration[4:0]) begin
            depthsOut_3 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h3 == iteration[4:0]) begin
              depthsOut_3 <= _GEN_66;
            end
          end else if (5'h3 == iteration[4:0]) begin
            depthsOut_3 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h4 == iteration[4:0]) begin
              depthsOut_4 <= 8'h20;
            end
          end else if (5'h4 == iteration[4:0]) begin
            depthsOut_4 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h4 == iteration[4:0]) begin
              depthsOut_4 <= _GEN_66;
            end
          end else if (5'h4 == iteration[4:0]) begin
            depthsOut_4 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h5 == iteration[4:0]) begin
              depthsOut_5 <= 8'h20;
            end
          end else if (5'h5 == iteration[4:0]) begin
            depthsOut_5 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h5 == iteration[4:0]) begin
              depthsOut_5 <= _GEN_66;
            end
          end else if (5'h5 == iteration[4:0]) begin
            depthsOut_5 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h6 == iteration[4:0]) begin
              depthsOut_6 <= 8'h20;
            end
          end else if (5'h6 == iteration[4:0]) begin
            depthsOut_6 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h6 == iteration[4:0]) begin
              depthsOut_6 <= _GEN_66;
            end
          end else if (5'h6 == iteration[4:0]) begin
            depthsOut_6 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h7 == iteration[4:0]) begin
              depthsOut_7 <= 8'h20;
            end
          end else if (5'h7 == iteration[4:0]) begin
            depthsOut_7 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h7 == iteration[4:0]) begin
              depthsOut_7 <= _GEN_66;
            end
          end else if (5'h7 == iteration[4:0]) begin
            depthsOut_7 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h8 == iteration[4:0]) begin
              depthsOut_8 <= 8'h20;
            end
          end else if (5'h8 == iteration[4:0]) begin
            depthsOut_8 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h8 == iteration[4:0]) begin
              depthsOut_8 <= _GEN_66;
            end
          end else if (5'h8 == iteration[4:0]) begin
            depthsOut_8 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h9 == iteration[4:0]) begin
              depthsOut_9 <= 8'h20;
            end
          end else if (5'h9 == iteration[4:0]) begin
            depthsOut_9 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h9 == iteration[4:0]) begin
              depthsOut_9 <= _GEN_66;
            end
          end else if (5'h9 == iteration[4:0]) begin
            depthsOut_9 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'ha == iteration[4:0]) begin
              depthsOut_10 <= 8'h20;
            end
          end else if (5'ha == iteration[4:0]) begin
            depthsOut_10 <= _GEN_66;
          end else if (_T_156) begin
            if (5'ha == iteration[4:0]) begin
              depthsOut_10 <= _GEN_66;
            end
          end else if (5'ha == iteration[4:0]) begin
            depthsOut_10 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'hb == iteration[4:0]) begin
              depthsOut_11 <= 8'h20;
            end
          end else if (5'hb == iteration[4:0]) begin
            depthsOut_11 <= _GEN_66;
          end else if (_T_156) begin
            if (5'hb == iteration[4:0]) begin
              depthsOut_11 <= _GEN_66;
            end
          end else if (5'hb == iteration[4:0]) begin
            depthsOut_11 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'hc == iteration[4:0]) begin
              depthsOut_12 <= 8'h20;
            end
          end else if (5'hc == iteration[4:0]) begin
            depthsOut_12 <= _GEN_66;
          end else if (_T_156) begin
            if (5'hc == iteration[4:0]) begin
              depthsOut_12 <= _GEN_66;
            end
          end else if (5'hc == iteration[4:0]) begin
            depthsOut_12 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'hd == iteration[4:0]) begin
              depthsOut_13 <= 8'h20;
            end
          end else if (5'hd == iteration[4:0]) begin
            depthsOut_13 <= _GEN_66;
          end else if (_T_156) begin
            if (5'hd == iteration[4:0]) begin
              depthsOut_13 <= _GEN_66;
            end
          end else if (5'hd == iteration[4:0]) begin
            depthsOut_13 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'he == iteration[4:0]) begin
              depthsOut_14 <= 8'h20;
            end
          end else if (5'he == iteration[4:0]) begin
            depthsOut_14 <= _GEN_66;
          end else if (_T_156) begin
            if (5'he == iteration[4:0]) begin
              depthsOut_14 <= _GEN_66;
            end
          end else if (5'he == iteration[4:0]) begin
            depthsOut_14 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'hf == iteration[4:0]) begin
              depthsOut_15 <= 8'h20;
            end
          end else if (5'hf == iteration[4:0]) begin
            depthsOut_15 <= _GEN_66;
          end else if (_T_156) begin
            if (5'hf == iteration[4:0]) begin
              depthsOut_15 <= _GEN_66;
            end
          end else if (5'hf == iteration[4:0]) begin
            depthsOut_15 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h10 == iteration[4:0]) begin
              depthsOut_16 <= 8'h20;
            end
          end else if (5'h10 == iteration[4:0]) begin
            depthsOut_16 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h10 == iteration[4:0]) begin
              depthsOut_16 <= _GEN_66;
            end
          end else if (5'h10 == iteration[4:0]) begin
            depthsOut_16 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h11 == iteration[4:0]) begin
              depthsOut_17 <= 8'h20;
            end
          end else if (5'h11 == iteration[4:0]) begin
            depthsOut_17 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h11 == iteration[4:0]) begin
              depthsOut_17 <= _GEN_66;
            end
          end else if (5'h11 == iteration[4:0]) begin
            depthsOut_17 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h12 == iteration[4:0]) begin
              depthsOut_18 <= 8'h20;
            end
          end else if (5'h12 == iteration[4:0]) begin
            depthsOut_18 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h12 == iteration[4:0]) begin
              depthsOut_18 <= _GEN_66;
            end
          end else if (5'h12 == iteration[4:0]) begin
            depthsOut_18 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h13 == iteration[4:0]) begin
              depthsOut_19 <= 8'h20;
            end
          end else if (5'h13 == iteration[4:0]) begin
            depthsOut_19 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h13 == iteration[4:0]) begin
              depthsOut_19 <= _GEN_66;
            end
          end else if (5'h13 == iteration[4:0]) begin
            depthsOut_19 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h14 == iteration[4:0]) begin
              depthsOut_20 <= 8'h20;
            end
          end else if (5'h14 == iteration[4:0]) begin
            depthsOut_20 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h14 == iteration[4:0]) begin
              depthsOut_20 <= _GEN_66;
            end
          end else if (5'h14 == iteration[4:0]) begin
            depthsOut_20 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h15 == iteration[4:0]) begin
              depthsOut_21 <= 8'h20;
            end
          end else if (5'h15 == iteration[4:0]) begin
            depthsOut_21 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h15 == iteration[4:0]) begin
              depthsOut_21 <= _GEN_66;
            end
          end else if (5'h15 == iteration[4:0]) begin
            depthsOut_21 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h16 == iteration[4:0]) begin
              depthsOut_22 <= 8'h20;
            end
          end else if (5'h16 == iteration[4:0]) begin
            depthsOut_22 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h16 == iteration[4:0]) begin
              depthsOut_22 <= _GEN_66;
            end
          end else if (5'h16 == iteration[4:0]) begin
            depthsOut_22 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h17 == iteration[4:0]) begin
              depthsOut_23 <= 8'h20;
            end
          end else if (5'h17 == iteration[4:0]) begin
            depthsOut_23 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h17 == iteration[4:0]) begin
              depthsOut_23 <= _GEN_66;
            end
          end else if (5'h17 == iteration[4:0]) begin
            depthsOut_23 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h18 == iteration[4:0]) begin
              depthsOut_24 <= 8'h20;
            end
          end else if (5'h18 == iteration[4:0]) begin
            depthsOut_24 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h18 == iteration[4:0]) begin
              depthsOut_24 <= _GEN_66;
            end
          end else if (5'h18 == iteration[4:0]) begin
            depthsOut_24 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h19 == iteration[4:0]) begin
              depthsOut_25 <= 8'h20;
            end
          end else if (5'h19 == iteration[4:0]) begin
            depthsOut_25 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h19 == iteration[4:0]) begin
              depthsOut_25 <= _GEN_66;
            end
          end else if (5'h19 == iteration[4:0]) begin
            depthsOut_25 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h1a == iteration[4:0]) begin
              depthsOut_26 <= 8'h20;
            end
          end else if (5'h1a == iteration[4:0]) begin
            depthsOut_26 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h1a == iteration[4:0]) begin
              depthsOut_26 <= _GEN_66;
            end
          end else if (5'h1a == iteration[4:0]) begin
            depthsOut_26 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h1b == iteration[4:0]) begin
              depthsOut_27 <= 8'h20;
            end
          end else if (5'h1b == iteration[4:0]) begin
            depthsOut_27 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h1b == iteration[4:0]) begin
              depthsOut_27 <= _GEN_66;
            end
          end else if (5'h1b == iteration[4:0]) begin
            depthsOut_27 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h1c == iteration[4:0]) begin
              depthsOut_28 <= 8'h20;
            end
          end else if (5'h1c == iteration[4:0]) begin
            depthsOut_28 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h1c == iteration[4:0]) begin
              depthsOut_28 <= _GEN_66;
            end
          end else if (5'h1c == iteration[4:0]) begin
            depthsOut_28 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h1d == iteration[4:0]) begin
              depthsOut_29 <= 8'h20;
            end
          end else if (5'h1d == iteration[4:0]) begin
            depthsOut_29 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h1d == iteration[4:0]) begin
              depthsOut_29 <= _GEN_66;
            end
          end else if (5'h1d == iteration[4:0]) begin
            depthsOut_29 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h1e == iteration[4:0]) begin
              depthsOut_30 <= 8'h20;
            end
          end else if (5'h1e == iteration[4:0]) begin
            depthsOut_30 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h1e == iteration[4:0]) begin
              depthsOut_30 <= _GEN_66;
            end
          end else if (5'h1e == iteration[4:0]) begin
            depthsOut_30 <= _T_162;
          end
        end
      end
    end
    if (!(_T_130)) begin
      if (!(_T_132)) begin
        if (_T_152) begin
          if (_T_134) begin
            if (5'h1f == iteration[4:0]) begin
              depthsOut_31 <= 8'h20;
            end
          end else if (5'h1f == iteration[4:0]) begin
            depthsOut_31 <= _GEN_66;
          end else if (_T_156) begin
            if (5'h1f == iteration[4:0]) begin
              depthsOut_31 <= _GEN_66;
            end
          end else if (5'h1f == iteration[4:0]) begin
            depthsOut_31 <= _T_162;
          end
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_0 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h0 == iteration[4:0]) begin
          charactersAtDepth_0 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_1 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h1 == iteration[4:0]) begin
          charactersAtDepth_1 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_2 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h2 == iteration[4:0]) begin
          charactersAtDepth_2 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_3 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h3 == iteration[4:0]) begin
          charactersAtDepth_3 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_4 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h4 == iteration[4:0]) begin
          charactersAtDepth_4 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_5 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h5 == iteration[4:0]) begin
          charactersAtDepth_5 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_6 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h6 == iteration[4:0]) begin
          charactersAtDepth_6 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_7 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h7 == iteration[4:0]) begin
          charactersAtDepth_7 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_8 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h8 == iteration[4:0]) begin
          charactersAtDepth_8 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_9 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h9 == iteration[4:0]) begin
          charactersAtDepth_9 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_10 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'ha == iteration[4:0]) begin
          charactersAtDepth_10 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_11 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'hb == iteration[4:0]) begin
          charactersAtDepth_11 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_12 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'hc == iteration[4:0]) begin
          charactersAtDepth_12 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_13 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'hd == iteration[4:0]) begin
          charactersAtDepth_13 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_14 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'he == iteration[4:0]) begin
          charactersAtDepth_14 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_15 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'hf == iteration[4:0]) begin
          charactersAtDepth_15 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_16 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h10 == iteration[4:0]) begin
          charactersAtDepth_16 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_17 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h11 == iteration[4:0]) begin
          charactersAtDepth_17 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_18 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h12 == iteration[4:0]) begin
          charactersAtDepth_18 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_19 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h13 == iteration[4:0]) begin
          charactersAtDepth_19 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_20 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h14 == iteration[4:0]) begin
          charactersAtDepth_20 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_21 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h15 == iteration[4:0]) begin
          charactersAtDepth_21 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_22 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h16 == iteration[4:0]) begin
          charactersAtDepth_22 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_23 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h17 == iteration[4:0]) begin
          charactersAtDepth_23 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_24 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h18 == iteration[4:0]) begin
          charactersAtDepth_24 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_25 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h19 == iteration[4:0]) begin
          charactersAtDepth_25 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_26 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h1a == iteration[4:0]) begin
          charactersAtDepth_26 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_27 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h1b == iteration[4:0]) begin
          charactersAtDepth_27 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_28 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h1c == iteration[4:0]) begin
          charactersAtDepth_28 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_29 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h1d == iteration[4:0]) begin
          charactersAtDepth_29 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_30 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (!(_T_134)) begin
        if (5'h1e == iteration[4:0]) begin
          charactersAtDepth_30 <= _T_142;
        end
      end
    end
    if (_T_130) begin
      if (io_start) begin
        charactersAtDepth_31 <= 6'sh0;
      end
    end else if (_T_132) begin
      if (_T_134) begin
        charactersAtDepth_31 <= _T_137;
      end else if (5'h1f == iteration[4:0]) begin
        charactersAtDepth_31 <= _T_142;
      end
    end
    if (_T_130) begin
      if (io_start) begin
        iteration <= 6'h0;
      end
    end else if (_T_132) begin
      if (!(_T_151)) begin
        iteration <= _T_144;
      end
    end else if (_T_152) begin
      iteration <= _T_166;
    end
  end
endmodule
module codewordGenerator(
  input         clock,
  input         reset,
  input         io_start,
  input  [8:0]  io_inputs_charactersOut_0,
  input  [8:0]  io_inputs_charactersOut_1,
  input  [8:0]  io_inputs_charactersOut_2,
  input  [8:0]  io_inputs_charactersOut_3,
  input  [8:0]  io_inputs_charactersOut_4,
  input  [8:0]  io_inputs_charactersOut_5,
  input  [8:0]  io_inputs_charactersOut_6,
  input  [8:0]  io_inputs_charactersOut_7,
  input  [8:0]  io_inputs_charactersOut_8,
  input  [8:0]  io_inputs_charactersOut_9,
  input  [8:0]  io_inputs_charactersOut_10,
  input  [8:0]  io_inputs_charactersOut_11,
  input  [8:0]  io_inputs_charactersOut_12,
  input  [8:0]  io_inputs_charactersOut_13,
  input  [8:0]  io_inputs_charactersOut_14,
  input  [8:0]  io_inputs_charactersOut_15,
  input  [8:0]  io_inputs_charactersOut_16,
  input  [8:0]  io_inputs_charactersOut_17,
  input  [8:0]  io_inputs_charactersOut_18,
  input  [8:0]  io_inputs_charactersOut_19,
  input  [8:0]  io_inputs_charactersOut_20,
  input  [8:0]  io_inputs_charactersOut_21,
  input  [8:0]  io_inputs_charactersOut_22,
  input  [8:0]  io_inputs_charactersOut_23,
  input  [8:0]  io_inputs_charactersOut_24,
  input  [8:0]  io_inputs_charactersOut_25,
  input  [8:0]  io_inputs_charactersOut_26,
  input  [8:0]  io_inputs_charactersOut_27,
  input  [8:0]  io_inputs_charactersOut_28,
  input  [8:0]  io_inputs_charactersOut_29,
  input  [8:0]  io_inputs_charactersOut_30,
  input  [8:0]  io_inputs_charactersOut_31,
  input  [7:0]  io_inputs_depthsOut_0,
  input  [7:0]  io_inputs_depthsOut_1,
  input  [7:0]  io_inputs_depthsOut_2,
  input  [7:0]  io_inputs_depthsOut_3,
  input  [7:0]  io_inputs_depthsOut_4,
  input  [7:0]  io_inputs_depthsOut_5,
  input  [7:0]  io_inputs_depthsOut_6,
  input  [7:0]  io_inputs_depthsOut_7,
  input  [7:0]  io_inputs_depthsOut_8,
  input  [7:0]  io_inputs_depthsOut_9,
  input  [7:0]  io_inputs_depthsOut_10,
  input  [7:0]  io_inputs_depthsOut_11,
  input  [7:0]  io_inputs_depthsOut_12,
  input  [7:0]  io_inputs_depthsOut_13,
  input  [7:0]  io_inputs_depthsOut_14,
  input  [7:0]  io_inputs_depthsOut_15,
  input  [7:0]  io_inputs_depthsOut_16,
  input  [7:0]  io_inputs_depthsOut_17,
  input  [7:0]  io_inputs_depthsOut_18,
  input  [7:0]  io_inputs_depthsOut_19,
  input  [7:0]  io_inputs_depthsOut_20,
  input  [7:0]  io_inputs_depthsOut_21,
  input  [7:0]  io_inputs_depthsOut_22,
  input  [7:0]  io_inputs_depthsOut_23,
  input  [7:0]  io_inputs_depthsOut_24,
  input  [7:0]  io_inputs_depthsOut_25,
  input  [7:0]  io_inputs_depthsOut_26,
  input  [7:0]  io_inputs_depthsOut_27,
  input  [7:0]  io_inputs_depthsOut_28,
  input  [7:0]  io_inputs_depthsOut_29,
  input  [7:0]  io_inputs_depthsOut_30,
  input  [7:0]  io_inputs_depthsOut_31,
  input  [8:0]  io_inputs_validNodesOut,
  output [23:0] io_outputs_codewords_0,
  output [23:0] io_outputs_codewords_1,
  output [23:0] io_outputs_codewords_2,
  output [23:0] io_outputs_codewords_3,
  output [23:0] io_outputs_codewords_4,
  output [23:0] io_outputs_codewords_5,
  output [23:0] io_outputs_codewords_6,
  output [23:0] io_outputs_codewords_7,
  output [23:0] io_outputs_codewords_8,
  output [23:0] io_outputs_codewords_9,
  output [23:0] io_outputs_codewords_10,
  output [23:0] io_outputs_codewords_11,
  output [23:0] io_outputs_codewords_12,
  output [23:0] io_outputs_codewords_13,
  output [23:0] io_outputs_codewords_14,
  output [23:0] io_outputs_codewords_15,
  output [23:0] io_outputs_codewords_16,
  output [23:0] io_outputs_codewords_17,
  output [23:0] io_outputs_codewords_18,
  output [23:0] io_outputs_codewords_19,
  output [23:0] io_outputs_codewords_20,
  output [23:0] io_outputs_codewords_21,
  output [23:0] io_outputs_codewords_22,
  output [23:0] io_outputs_codewords_23,
  output [23:0] io_outputs_codewords_24,
  output [23:0] io_outputs_codewords_25,
  output [23:0] io_outputs_codewords_26,
  output [23:0] io_outputs_codewords_27,
  output [23:0] io_outputs_codewords_28,
  output [23:0] io_outputs_codewords_29,
  output [23:0] io_outputs_codewords_30,
  output [23:0] io_outputs_codewords_31,
  output [23:0] io_outputs_codewords_32,
  output [23:0] io_outputs_codewords_33,
  output [23:0] io_outputs_codewords_34,
  output [23:0] io_outputs_codewords_35,
  output [23:0] io_outputs_codewords_36,
  output [23:0] io_outputs_codewords_37,
  output [23:0] io_outputs_codewords_38,
  output [23:0] io_outputs_codewords_39,
  output [23:0] io_outputs_codewords_40,
  output [23:0] io_outputs_codewords_41,
  output [23:0] io_outputs_codewords_42,
  output [23:0] io_outputs_codewords_43,
  output [23:0] io_outputs_codewords_44,
  output [23:0] io_outputs_codewords_45,
  output [23:0] io_outputs_codewords_46,
  output [23:0] io_outputs_codewords_47,
  output [23:0] io_outputs_codewords_48,
  output [23:0] io_outputs_codewords_49,
  output [23:0] io_outputs_codewords_50,
  output [23:0] io_outputs_codewords_51,
  output [23:0] io_outputs_codewords_52,
  output [23:0] io_outputs_codewords_53,
  output [23:0] io_outputs_codewords_54,
  output [23:0] io_outputs_codewords_55,
  output [23:0] io_outputs_codewords_56,
  output [23:0] io_outputs_codewords_57,
  output [23:0] io_outputs_codewords_58,
  output [23:0] io_outputs_codewords_59,
  output [23:0] io_outputs_codewords_60,
  output [23:0] io_outputs_codewords_61,
  output [23:0] io_outputs_codewords_62,
  output [23:0] io_outputs_codewords_63,
  output [23:0] io_outputs_codewords_64,
  output [23:0] io_outputs_codewords_65,
  output [23:0] io_outputs_codewords_66,
  output [23:0] io_outputs_codewords_67,
  output [23:0] io_outputs_codewords_68,
  output [23:0] io_outputs_codewords_69,
  output [23:0] io_outputs_codewords_70,
  output [23:0] io_outputs_codewords_71,
  output [23:0] io_outputs_codewords_72,
  output [23:0] io_outputs_codewords_73,
  output [23:0] io_outputs_codewords_74,
  output [23:0] io_outputs_codewords_75,
  output [23:0] io_outputs_codewords_76,
  output [23:0] io_outputs_codewords_77,
  output [23:0] io_outputs_codewords_78,
  output [23:0] io_outputs_codewords_79,
  output [23:0] io_outputs_codewords_80,
  output [23:0] io_outputs_codewords_81,
  output [23:0] io_outputs_codewords_82,
  output [23:0] io_outputs_codewords_83,
  output [23:0] io_outputs_codewords_84,
  output [23:0] io_outputs_codewords_85,
  output [23:0] io_outputs_codewords_86,
  output [23:0] io_outputs_codewords_87,
  output [23:0] io_outputs_codewords_88,
  output [23:0] io_outputs_codewords_89,
  output [23:0] io_outputs_codewords_90,
  output [23:0] io_outputs_codewords_91,
  output [23:0] io_outputs_codewords_92,
  output [23:0] io_outputs_codewords_93,
  output [23:0] io_outputs_codewords_94,
  output [23:0] io_outputs_codewords_95,
  output [23:0] io_outputs_codewords_96,
  output [23:0] io_outputs_codewords_97,
  output [23:0] io_outputs_codewords_98,
  output [23:0] io_outputs_codewords_99,
  output [23:0] io_outputs_codewords_100,
  output [23:0] io_outputs_codewords_101,
  output [23:0] io_outputs_codewords_102,
  output [23:0] io_outputs_codewords_103,
  output [23:0] io_outputs_codewords_104,
  output [23:0] io_outputs_codewords_105,
  output [23:0] io_outputs_codewords_106,
  output [23:0] io_outputs_codewords_107,
  output [23:0] io_outputs_codewords_108,
  output [23:0] io_outputs_codewords_109,
  output [23:0] io_outputs_codewords_110,
  output [23:0] io_outputs_codewords_111,
  output [23:0] io_outputs_codewords_112,
  output [23:0] io_outputs_codewords_113,
  output [23:0] io_outputs_codewords_114,
  output [23:0] io_outputs_codewords_115,
  output [23:0] io_outputs_codewords_116,
  output [23:0] io_outputs_codewords_117,
  output [23:0] io_outputs_codewords_118,
  output [23:0] io_outputs_codewords_119,
  output [23:0] io_outputs_codewords_120,
  output [23:0] io_outputs_codewords_121,
  output [23:0] io_outputs_codewords_122,
  output [23:0] io_outputs_codewords_123,
  output [23:0] io_outputs_codewords_124,
  output [23:0] io_outputs_codewords_125,
  output [23:0] io_outputs_codewords_126,
  output [23:0] io_outputs_codewords_127,
  output [23:0] io_outputs_codewords_128,
  output [23:0] io_outputs_codewords_129,
  output [23:0] io_outputs_codewords_130,
  output [23:0] io_outputs_codewords_131,
  output [23:0] io_outputs_codewords_132,
  output [23:0] io_outputs_codewords_133,
  output [23:0] io_outputs_codewords_134,
  output [23:0] io_outputs_codewords_135,
  output [23:0] io_outputs_codewords_136,
  output [23:0] io_outputs_codewords_137,
  output [23:0] io_outputs_codewords_138,
  output [23:0] io_outputs_codewords_139,
  output [23:0] io_outputs_codewords_140,
  output [23:0] io_outputs_codewords_141,
  output [23:0] io_outputs_codewords_142,
  output [23:0] io_outputs_codewords_143,
  output [23:0] io_outputs_codewords_144,
  output [23:0] io_outputs_codewords_145,
  output [23:0] io_outputs_codewords_146,
  output [23:0] io_outputs_codewords_147,
  output [23:0] io_outputs_codewords_148,
  output [23:0] io_outputs_codewords_149,
  output [23:0] io_outputs_codewords_150,
  output [23:0] io_outputs_codewords_151,
  output [23:0] io_outputs_codewords_152,
  output [23:0] io_outputs_codewords_153,
  output [23:0] io_outputs_codewords_154,
  output [23:0] io_outputs_codewords_155,
  output [23:0] io_outputs_codewords_156,
  output [23:0] io_outputs_codewords_157,
  output [23:0] io_outputs_codewords_158,
  output [23:0] io_outputs_codewords_159,
  output [23:0] io_outputs_codewords_160,
  output [23:0] io_outputs_codewords_161,
  output [23:0] io_outputs_codewords_162,
  output [23:0] io_outputs_codewords_163,
  output [23:0] io_outputs_codewords_164,
  output [23:0] io_outputs_codewords_165,
  output [23:0] io_outputs_codewords_166,
  output [23:0] io_outputs_codewords_167,
  output [23:0] io_outputs_codewords_168,
  output [23:0] io_outputs_codewords_169,
  output [23:0] io_outputs_codewords_170,
  output [23:0] io_outputs_codewords_171,
  output [23:0] io_outputs_codewords_172,
  output [23:0] io_outputs_codewords_173,
  output [23:0] io_outputs_codewords_174,
  output [23:0] io_outputs_codewords_175,
  output [23:0] io_outputs_codewords_176,
  output [23:0] io_outputs_codewords_177,
  output [23:0] io_outputs_codewords_178,
  output [23:0] io_outputs_codewords_179,
  output [23:0] io_outputs_codewords_180,
  output [23:0] io_outputs_codewords_181,
  output [23:0] io_outputs_codewords_182,
  output [23:0] io_outputs_codewords_183,
  output [23:0] io_outputs_codewords_184,
  output [23:0] io_outputs_codewords_185,
  output [23:0] io_outputs_codewords_186,
  output [23:0] io_outputs_codewords_187,
  output [23:0] io_outputs_codewords_188,
  output [23:0] io_outputs_codewords_189,
  output [23:0] io_outputs_codewords_190,
  output [23:0] io_outputs_codewords_191,
  output [23:0] io_outputs_codewords_192,
  output [23:0] io_outputs_codewords_193,
  output [23:0] io_outputs_codewords_194,
  output [23:0] io_outputs_codewords_195,
  output [23:0] io_outputs_codewords_196,
  output [23:0] io_outputs_codewords_197,
  output [23:0] io_outputs_codewords_198,
  output [23:0] io_outputs_codewords_199,
  output [23:0] io_outputs_codewords_200,
  output [23:0] io_outputs_codewords_201,
  output [23:0] io_outputs_codewords_202,
  output [23:0] io_outputs_codewords_203,
  output [23:0] io_outputs_codewords_204,
  output [23:0] io_outputs_codewords_205,
  output [23:0] io_outputs_codewords_206,
  output [23:0] io_outputs_codewords_207,
  output [23:0] io_outputs_codewords_208,
  output [23:0] io_outputs_codewords_209,
  output [23:0] io_outputs_codewords_210,
  output [23:0] io_outputs_codewords_211,
  output [23:0] io_outputs_codewords_212,
  output [23:0] io_outputs_codewords_213,
  output [23:0] io_outputs_codewords_214,
  output [23:0] io_outputs_codewords_215,
  output [23:0] io_outputs_codewords_216,
  output [23:0] io_outputs_codewords_217,
  output [23:0] io_outputs_codewords_218,
  output [23:0] io_outputs_codewords_219,
  output [23:0] io_outputs_codewords_220,
  output [23:0] io_outputs_codewords_221,
  output [23:0] io_outputs_codewords_222,
  output [23:0] io_outputs_codewords_223,
  output [23:0] io_outputs_codewords_224,
  output [23:0] io_outputs_codewords_225,
  output [23:0] io_outputs_codewords_226,
  output [23:0] io_outputs_codewords_227,
  output [23:0] io_outputs_codewords_228,
  output [23:0] io_outputs_codewords_229,
  output [23:0] io_outputs_codewords_230,
  output [23:0] io_outputs_codewords_231,
  output [23:0] io_outputs_codewords_232,
  output [23:0] io_outputs_codewords_233,
  output [23:0] io_outputs_codewords_234,
  output [23:0] io_outputs_codewords_235,
  output [23:0] io_outputs_codewords_236,
  output [23:0] io_outputs_codewords_237,
  output [23:0] io_outputs_codewords_238,
  output [23:0] io_outputs_codewords_239,
  output [23:0] io_outputs_codewords_240,
  output [23:0] io_outputs_codewords_241,
  output [23:0] io_outputs_codewords_242,
  output [23:0] io_outputs_codewords_243,
  output [23:0] io_outputs_codewords_244,
  output [23:0] io_outputs_codewords_245,
  output [23:0] io_outputs_codewords_246,
  output [23:0] io_outputs_codewords_247,
  output [23:0] io_outputs_codewords_248,
  output [23:0] io_outputs_codewords_249,
  output [23:0] io_outputs_codewords_250,
  output [23:0] io_outputs_codewords_251,
  output [23:0] io_outputs_codewords_252,
  output [23:0] io_outputs_codewords_253,
  output [23:0] io_outputs_codewords_254,
  output [23:0] io_outputs_codewords_255,
  output [4:0]  io_outputs_lengths_0,
  output [4:0]  io_outputs_lengths_1,
  output [4:0]  io_outputs_lengths_2,
  output [4:0]  io_outputs_lengths_3,
  output [4:0]  io_outputs_lengths_4,
  output [4:0]  io_outputs_lengths_5,
  output [4:0]  io_outputs_lengths_6,
  output [4:0]  io_outputs_lengths_7,
  output [4:0]  io_outputs_lengths_8,
  output [4:0]  io_outputs_lengths_9,
  output [4:0]  io_outputs_lengths_10,
  output [4:0]  io_outputs_lengths_11,
  output [4:0]  io_outputs_lengths_12,
  output [4:0]  io_outputs_lengths_13,
  output [4:0]  io_outputs_lengths_14,
  output [4:0]  io_outputs_lengths_15,
  output [4:0]  io_outputs_lengths_16,
  output [4:0]  io_outputs_lengths_17,
  output [4:0]  io_outputs_lengths_18,
  output [4:0]  io_outputs_lengths_19,
  output [4:0]  io_outputs_lengths_20,
  output [4:0]  io_outputs_lengths_21,
  output [4:0]  io_outputs_lengths_22,
  output [4:0]  io_outputs_lengths_23,
  output [4:0]  io_outputs_lengths_24,
  output [4:0]  io_outputs_lengths_25,
  output [4:0]  io_outputs_lengths_26,
  output [4:0]  io_outputs_lengths_27,
  output [4:0]  io_outputs_lengths_28,
  output [4:0]  io_outputs_lengths_29,
  output [4:0]  io_outputs_lengths_30,
  output [4:0]  io_outputs_lengths_31,
  output [4:0]  io_outputs_lengths_32,
  output [4:0]  io_outputs_lengths_33,
  output [4:0]  io_outputs_lengths_34,
  output [4:0]  io_outputs_lengths_35,
  output [4:0]  io_outputs_lengths_36,
  output [4:0]  io_outputs_lengths_37,
  output [4:0]  io_outputs_lengths_38,
  output [4:0]  io_outputs_lengths_39,
  output [4:0]  io_outputs_lengths_40,
  output [4:0]  io_outputs_lengths_41,
  output [4:0]  io_outputs_lengths_42,
  output [4:0]  io_outputs_lengths_43,
  output [4:0]  io_outputs_lengths_44,
  output [4:0]  io_outputs_lengths_45,
  output [4:0]  io_outputs_lengths_46,
  output [4:0]  io_outputs_lengths_47,
  output [4:0]  io_outputs_lengths_48,
  output [4:0]  io_outputs_lengths_49,
  output [4:0]  io_outputs_lengths_50,
  output [4:0]  io_outputs_lengths_51,
  output [4:0]  io_outputs_lengths_52,
  output [4:0]  io_outputs_lengths_53,
  output [4:0]  io_outputs_lengths_54,
  output [4:0]  io_outputs_lengths_55,
  output [4:0]  io_outputs_lengths_56,
  output [4:0]  io_outputs_lengths_57,
  output [4:0]  io_outputs_lengths_58,
  output [4:0]  io_outputs_lengths_59,
  output [4:0]  io_outputs_lengths_60,
  output [4:0]  io_outputs_lengths_61,
  output [4:0]  io_outputs_lengths_62,
  output [4:0]  io_outputs_lengths_63,
  output [4:0]  io_outputs_lengths_64,
  output [4:0]  io_outputs_lengths_65,
  output [4:0]  io_outputs_lengths_66,
  output [4:0]  io_outputs_lengths_67,
  output [4:0]  io_outputs_lengths_68,
  output [4:0]  io_outputs_lengths_69,
  output [4:0]  io_outputs_lengths_70,
  output [4:0]  io_outputs_lengths_71,
  output [4:0]  io_outputs_lengths_72,
  output [4:0]  io_outputs_lengths_73,
  output [4:0]  io_outputs_lengths_74,
  output [4:0]  io_outputs_lengths_75,
  output [4:0]  io_outputs_lengths_76,
  output [4:0]  io_outputs_lengths_77,
  output [4:0]  io_outputs_lengths_78,
  output [4:0]  io_outputs_lengths_79,
  output [4:0]  io_outputs_lengths_80,
  output [4:0]  io_outputs_lengths_81,
  output [4:0]  io_outputs_lengths_82,
  output [4:0]  io_outputs_lengths_83,
  output [4:0]  io_outputs_lengths_84,
  output [4:0]  io_outputs_lengths_85,
  output [4:0]  io_outputs_lengths_86,
  output [4:0]  io_outputs_lengths_87,
  output [4:0]  io_outputs_lengths_88,
  output [4:0]  io_outputs_lengths_89,
  output [4:0]  io_outputs_lengths_90,
  output [4:0]  io_outputs_lengths_91,
  output [4:0]  io_outputs_lengths_92,
  output [4:0]  io_outputs_lengths_93,
  output [4:0]  io_outputs_lengths_94,
  output [4:0]  io_outputs_lengths_95,
  output [4:0]  io_outputs_lengths_96,
  output [4:0]  io_outputs_lengths_97,
  output [4:0]  io_outputs_lengths_98,
  output [4:0]  io_outputs_lengths_99,
  output [4:0]  io_outputs_lengths_100,
  output [4:0]  io_outputs_lengths_101,
  output [4:0]  io_outputs_lengths_102,
  output [4:0]  io_outputs_lengths_103,
  output [4:0]  io_outputs_lengths_104,
  output [4:0]  io_outputs_lengths_105,
  output [4:0]  io_outputs_lengths_106,
  output [4:0]  io_outputs_lengths_107,
  output [4:0]  io_outputs_lengths_108,
  output [4:0]  io_outputs_lengths_109,
  output [4:0]  io_outputs_lengths_110,
  output [4:0]  io_outputs_lengths_111,
  output [4:0]  io_outputs_lengths_112,
  output [4:0]  io_outputs_lengths_113,
  output [4:0]  io_outputs_lengths_114,
  output [4:0]  io_outputs_lengths_115,
  output [4:0]  io_outputs_lengths_116,
  output [4:0]  io_outputs_lengths_117,
  output [4:0]  io_outputs_lengths_118,
  output [4:0]  io_outputs_lengths_119,
  output [4:0]  io_outputs_lengths_120,
  output [4:0]  io_outputs_lengths_121,
  output [4:0]  io_outputs_lengths_122,
  output [4:0]  io_outputs_lengths_123,
  output [4:0]  io_outputs_lengths_124,
  output [4:0]  io_outputs_lengths_125,
  output [4:0]  io_outputs_lengths_126,
  output [4:0]  io_outputs_lengths_127,
  output [4:0]  io_outputs_lengths_128,
  output [4:0]  io_outputs_lengths_129,
  output [4:0]  io_outputs_lengths_130,
  output [4:0]  io_outputs_lengths_131,
  output [4:0]  io_outputs_lengths_132,
  output [4:0]  io_outputs_lengths_133,
  output [4:0]  io_outputs_lengths_134,
  output [4:0]  io_outputs_lengths_135,
  output [4:0]  io_outputs_lengths_136,
  output [4:0]  io_outputs_lengths_137,
  output [4:0]  io_outputs_lengths_138,
  output [4:0]  io_outputs_lengths_139,
  output [4:0]  io_outputs_lengths_140,
  output [4:0]  io_outputs_lengths_141,
  output [4:0]  io_outputs_lengths_142,
  output [4:0]  io_outputs_lengths_143,
  output [4:0]  io_outputs_lengths_144,
  output [4:0]  io_outputs_lengths_145,
  output [4:0]  io_outputs_lengths_146,
  output [4:0]  io_outputs_lengths_147,
  output [4:0]  io_outputs_lengths_148,
  output [4:0]  io_outputs_lengths_149,
  output [4:0]  io_outputs_lengths_150,
  output [4:0]  io_outputs_lengths_151,
  output [4:0]  io_outputs_lengths_152,
  output [4:0]  io_outputs_lengths_153,
  output [4:0]  io_outputs_lengths_154,
  output [4:0]  io_outputs_lengths_155,
  output [4:0]  io_outputs_lengths_156,
  output [4:0]  io_outputs_lengths_157,
  output [4:0]  io_outputs_lengths_158,
  output [4:0]  io_outputs_lengths_159,
  output [4:0]  io_outputs_lengths_160,
  output [4:0]  io_outputs_lengths_161,
  output [4:0]  io_outputs_lengths_162,
  output [4:0]  io_outputs_lengths_163,
  output [4:0]  io_outputs_lengths_164,
  output [4:0]  io_outputs_lengths_165,
  output [4:0]  io_outputs_lengths_166,
  output [4:0]  io_outputs_lengths_167,
  output [4:0]  io_outputs_lengths_168,
  output [4:0]  io_outputs_lengths_169,
  output [4:0]  io_outputs_lengths_170,
  output [4:0]  io_outputs_lengths_171,
  output [4:0]  io_outputs_lengths_172,
  output [4:0]  io_outputs_lengths_173,
  output [4:0]  io_outputs_lengths_174,
  output [4:0]  io_outputs_lengths_175,
  output [4:0]  io_outputs_lengths_176,
  output [4:0]  io_outputs_lengths_177,
  output [4:0]  io_outputs_lengths_178,
  output [4:0]  io_outputs_lengths_179,
  output [4:0]  io_outputs_lengths_180,
  output [4:0]  io_outputs_lengths_181,
  output [4:0]  io_outputs_lengths_182,
  output [4:0]  io_outputs_lengths_183,
  output [4:0]  io_outputs_lengths_184,
  output [4:0]  io_outputs_lengths_185,
  output [4:0]  io_outputs_lengths_186,
  output [4:0]  io_outputs_lengths_187,
  output [4:0]  io_outputs_lengths_188,
  output [4:0]  io_outputs_lengths_189,
  output [4:0]  io_outputs_lengths_190,
  output [4:0]  io_outputs_lengths_191,
  output [4:0]  io_outputs_lengths_192,
  output [4:0]  io_outputs_lengths_193,
  output [4:0]  io_outputs_lengths_194,
  output [4:0]  io_outputs_lengths_195,
  output [4:0]  io_outputs_lengths_196,
  output [4:0]  io_outputs_lengths_197,
  output [4:0]  io_outputs_lengths_198,
  output [4:0]  io_outputs_lengths_199,
  output [4:0]  io_outputs_lengths_200,
  output [4:0]  io_outputs_lengths_201,
  output [4:0]  io_outputs_lengths_202,
  output [4:0]  io_outputs_lengths_203,
  output [4:0]  io_outputs_lengths_204,
  output [4:0]  io_outputs_lengths_205,
  output [4:0]  io_outputs_lengths_206,
  output [4:0]  io_outputs_lengths_207,
  output [4:0]  io_outputs_lengths_208,
  output [4:0]  io_outputs_lengths_209,
  output [4:0]  io_outputs_lengths_210,
  output [4:0]  io_outputs_lengths_211,
  output [4:0]  io_outputs_lengths_212,
  output [4:0]  io_outputs_lengths_213,
  output [4:0]  io_outputs_lengths_214,
  output [4:0]  io_outputs_lengths_215,
  output [4:0]  io_outputs_lengths_216,
  output [4:0]  io_outputs_lengths_217,
  output [4:0]  io_outputs_lengths_218,
  output [4:0]  io_outputs_lengths_219,
  output [4:0]  io_outputs_lengths_220,
  output [4:0]  io_outputs_lengths_221,
  output [4:0]  io_outputs_lengths_222,
  output [4:0]  io_outputs_lengths_223,
  output [4:0]  io_outputs_lengths_224,
  output [4:0]  io_outputs_lengths_225,
  output [4:0]  io_outputs_lengths_226,
  output [4:0]  io_outputs_lengths_227,
  output [4:0]  io_outputs_lengths_228,
  output [4:0]  io_outputs_lengths_229,
  output [4:0]  io_outputs_lengths_230,
  output [4:0]  io_outputs_lengths_231,
  output [4:0]  io_outputs_lengths_232,
  output [4:0]  io_outputs_lengths_233,
  output [4:0]  io_outputs_lengths_234,
  output [4:0]  io_outputs_lengths_235,
  output [4:0]  io_outputs_lengths_236,
  output [4:0]  io_outputs_lengths_237,
  output [4:0]  io_outputs_lengths_238,
  output [4:0]  io_outputs_lengths_239,
  output [4:0]  io_outputs_lengths_240,
  output [4:0]  io_outputs_lengths_241,
  output [4:0]  io_outputs_lengths_242,
  output [4:0]  io_outputs_lengths_243,
  output [4:0]  io_outputs_lengths_244,
  output [4:0]  io_outputs_lengths_245,
  output [4:0]  io_outputs_lengths_246,
  output [4:0]  io_outputs_lengths_247,
  output [4:0]  io_outputs_lengths_248,
  output [4:0]  io_outputs_lengths_249,
  output [4:0]  io_outputs_lengths_250,
  output [4:0]  io_outputs_lengths_251,
  output [4:0]  io_outputs_lengths_252,
  output [4:0]  io_outputs_lengths_253,
  output [4:0]  io_outputs_lengths_254,
  output [4:0]  io_outputs_lengths_255,
  output [8:0]  io_outputs_charactersOut_0,
  output [8:0]  io_outputs_charactersOut_1,
  output [8:0]  io_outputs_charactersOut_2,
  output [8:0]  io_outputs_charactersOut_3,
  output [8:0]  io_outputs_charactersOut_4,
  output [8:0]  io_outputs_charactersOut_5,
  output [8:0]  io_outputs_charactersOut_6,
  output [8:0]  io_outputs_charactersOut_7,
  output [8:0]  io_outputs_charactersOut_8,
  output [8:0]  io_outputs_charactersOut_9,
  output [8:0]  io_outputs_charactersOut_10,
  output [8:0]  io_outputs_charactersOut_11,
  output [8:0]  io_outputs_charactersOut_12,
  output [8:0]  io_outputs_charactersOut_13,
  output [8:0]  io_outputs_charactersOut_14,
  output [8:0]  io_outputs_charactersOut_15,
  output [8:0]  io_outputs_charactersOut_16,
  output [8:0]  io_outputs_charactersOut_17,
  output [8:0]  io_outputs_charactersOut_18,
  output [8:0]  io_outputs_charactersOut_19,
  output [8:0]  io_outputs_charactersOut_20,
  output [8:0]  io_outputs_charactersOut_21,
  output [8:0]  io_outputs_charactersOut_22,
  output [8:0]  io_outputs_charactersOut_23,
  output [8:0]  io_outputs_charactersOut_24,
  output [8:0]  io_outputs_charactersOut_25,
  output [8:0]  io_outputs_charactersOut_26,
  output [8:0]  io_outputs_charactersOut_27,
  output [8:0]  io_outputs_charactersOut_28,
  output [8:0]  io_outputs_charactersOut_29,
  output [8:0]  io_outputs_charactersOut_30,
  output [8:0]  io_outputs_charactersOut_31,
  output [8:0]  io_outputs_nodes,
  output [3:0]  io_outputs_escapeCharacterLength,
  output [15:0] io_outputs_escapeCodeword,
  output        io_finished
);
  reg [1:0] state; // @[codewordGenerator.scala 37:22]
  reg [31:0] _RAND_0;
  reg [8:0] charactersIn_0; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_1;
  reg [8:0] charactersIn_1; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_2;
  reg [8:0] charactersIn_2; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_3;
  reg [8:0] charactersIn_3; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_4;
  reg [8:0] charactersIn_4; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_5;
  reg [8:0] charactersIn_5; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_6;
  reg [8:0] charactersIn_6; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_7;
  reg [8:0] charactersIn_7; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_8;
  reg [8:0] charactersIn_8; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_9;
  reg [8:0] charactersIn_9; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_10;
  reg [8:0] charactersIn_10; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_11;
  reg [8:0] charactersIn_11; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_12;
  reg [8:0] charactersIn_12; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_13;
  reg [8:0] charactersIn_13; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_14;
  reg [8:0] charactersIn_14; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_15;
  reg [8:0] charactersIn_15; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_16;
  reg [8:0] charactersIn_16; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_17;
  reg [8:0] charactersIn_17; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_18;
  reg [8:0] charactersIn_18; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_19;
  reg [8:0] charactersIn_19; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_20;
  reg [8:0] charactersIn_20; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_21;
  reg [8:0] charactersIn_21; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_22;
  reg [8:0] charactersIn_22; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_23;
  reg [8:0] charactersIn_23; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_24;
  reg [8:0] charactersIn_24; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_25;
  reg [8:0] charactersIn_25; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_26;
  reg [8:0] charactersIn_26; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_27;
  reg [8:0] charactersIn_27; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_28;
  reg [8:0] charactersIn_28; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_29;
  reg [8:0] charactersIn_29; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_30;
  reg [8:0] charactersIn_30; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_31;
  reg [8:0] charactersIn_31; // @[codewordGenerator.scala 40:29]
  reg [31:0] _RAND_32;
  reg [3:0] depths_0; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_33;
  reg [3:0] depths_1; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_34;
  reg [3:0] depths_2; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_35;
  reg [3:0] depths_3; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_36;
  reg [3:0] depths_4; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_37;
  reg [3:0] depths_5; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_38;
  reg [3:0] depths_6; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_39;
  reg [3:0] depths_7; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_40;
  reg [3:0] depths_8; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_41;
  reg [3:0] depths_9; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_42;
  reg [3:0] depths_10; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_43;
  reg [3:0] depths_11; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_44;
  reg [3:0] depths_12; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_45;
  reg [3:0] depths_13; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_46;
  reg [3:0] depths_14; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_47;
  reg [3:0] depths_15; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_48;
  reg [3:0] depths_16; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_49;
  reg [3:0] depths_17; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_50;
  reg [3:0] depths_18; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_51;
  reg [3:0] depths_19; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_52;
  reg [3:0] depths_20; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_53;
  reg [3:0] depths_21; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_54;
  reg [3:0] depths_22; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_55;
  reg [3:0] depths_23; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_56;
  reg [3:0] depths_24; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_57;
  reg [3:0] depths_25; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_58;
  reg [3:0] depths_26; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_59;
  reg [3:0] depths_27; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_60;
  reg [3:0] depths_28; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_61;
  reg [3:0] depths_29; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_62;
  reg [3:0] depths_30; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_63;
  reg [3:0] depths_31; // @[codewordGenerator.scala 45:23]
  reg [31:0] _RAND_64;
  reg [15:0] codewords_0; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_65;
  reg [15:0] codewords_1; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_66;
  reg [15:0] codewords_2; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_67;
  reg [15:0] codewords_3; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_68;
  reg [15:0] codewords_4; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_69;
  reg [15:0] codewords_5; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_70;
  reg [15:0] codewords_6; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_71;
  reg [15:0] codewords_7; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_72;
  reg [15:0] codewords_8; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_73;
  reg [15:0] codewords_9; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_74;
  reg [15:0] codewords_10; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_75;
  reg [15:0] codewords_11; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_76;
  reg [15:0] codewords_12; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_77;
  reg [15:0] codewords_13; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_78;
  reg [15:0] codewords_14; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_79;
  reg [15:0] codewords_15; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_80;
  reg [15:0] codewords_16; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_81;
  reg [15:0] codewords_17; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_82;
  reg [15:0] codewords_18; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_83;
  reg [15:0] codewords_19; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_84;
  reg [15:0] codewords_20; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_85;
  reg [15:0] codewords_21; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_86;
  reg [15:0] codewords_22; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_87;
  reg [15:0] codewords_23; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_88;
  reg [15:0] codewords_24; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_89;
  reg [15:0] codewords_25; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_90;
  reg [15:0] codewords_26; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_91;
  reg [15:0] codewords_27; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_92;
  reg [15:0] codewords_28; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_93;
  reg [15:0] codewords_29; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_94;
  reg [15:0] codewords_30; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_95;
  reg [15:0] codewords_31; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_96;
  reg [15:0] codewords_32; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_97;
  reg [15:0] codewords_33; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_98;
  reg [15:0] codewords_34; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_99;
  reg [15:0] codewords_35; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_100;
  reg [15:0] codewords_36; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_101;
  reg [15:0] codewords_37; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_102;
  reg [15:0] codewords_38; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_103;
  reg [15:0] codewords_39; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_104;
  reg [15:0] codewords_40; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_105;
  reg [15:0] codewords_41; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_106;
  reg [15:0] codewords_42; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_107;
  reg [15:0] codewords_43; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_108;
  reg [15:0] codewords_44; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_109;
  reg [15:0] codewords_45; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_110;
  reg [15:0] codewords_46; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_111;
  reg [15:0] codewords_47; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_112;
  reg [15:0] codewords_48; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_113;
  reg [15:0] codewords_49; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_114;
  reg [15:0] codewords_50; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_115;
  reg [15:0] codewords_51; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_116;
  reg [15:0] codewords_52; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_117;
  reg [15:0] codewords_53; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_118;
  reg [15:0] codewords_54; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_119;
  reg [15:0] codewords_55; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_120;
  reg [15:0] codewords_56; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_121;
  reg [15:0] codewords_57; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_122;
  reg [15:0] codewords_58; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_123;
  reg [15:0] codewords_59; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_124;
  reg [15:0] codewords_60; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_125;
  reg [15:0] codewords_61; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_126;
  reg [15:0] codewords_62; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_127;
  reg [15:0] codewords_63; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_128;
  reg [15:0] codewords_64; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_129;
  reg [15:0] codewords_65; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_130;
  reg [15:0] codewords_66; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_131;
  reg [15:0] codewords_67; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_132;
  reg [15:0] codewords_68; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_133;
  reg [15:0] codewords_69; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_134;
  reg [15:0] codewords_70; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_135;
  reg [15:0] codewords_71; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_136;
  reg [15:0] codewords_72; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_137;
  reg [15:0] codewords_73; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_138;
  reg [15:0] codewords_74; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_139;
  reg [15:0] codewords_75; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_140;
  reg [15:0] codewords_76; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_141;
  reg [15:0] codewords_77; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_142;
  reg [15:0] codewords_78; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_143;
  reg [15:0] codewords_79; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_144;
  reg [15:0] codewords_80; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_145;
  reg [15:0] codewords_81; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_146;
  reg [15:0] codewords_82; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_147;
  reg [15:0] codewords_83; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_148;
  reg [15:0] codewords_84; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_149;
  reg [15:0] codewords_85; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_150;
  reg [15:0] codewords_86; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_151;
  reg [15:0] codewords_87; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_152;
  reg [15:0] codewords_88; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_153;
  reg [15:0] codewords_89; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_154;
  reg [15:0] codewords_90; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_155;
  reg [15:0] codewords_91; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_156;
  reg [15:0] codewords_92; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_157;
  reg [15:0] codewords_93; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_158;
  reg [15:0] codewords_94; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_159;
  reg [15:0] codewords_95; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_160;
  reg [15:0] codewords_96; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_161;
  reg [15:0] codewords_97; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_162;
  reg [15:0] codewords_98; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_163;
  reg [15:0] codewords_99; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_164;
  reg [15:0] codewords_100; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_165;
  reg [15:0] codewords_101; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_166;
  reg [15:0] codewords_102; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_167;
  reg [15:0] codewords_103; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_168;
  reg [15:0] codewords_104; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_169;
  reg [15:0] codewords_105; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_170;
  reg [15:0] codewords_106; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_171;
  reg [15:0] codewords_107; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_172;
  reg [15:0] codewords_108; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_173;
  reg [15:0] codewords_109; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_174;
  reg [15:0] codewords_110; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_175;
  reg [15:0] codewords_111; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_176;
  reg [15:0] codewords_112; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_177;
  reg [15:0] codewords_113; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_178;
  reg [15:0] codewords_114; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_179;
  reg [15:0] codewords_115; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_180;
  reg [15:0] codewords_116; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_181;
  reg [15:0] codewords_117; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_182;
  reg [15:0] codewords_118; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_183;
  reg [15:0] codewords_119; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_184;
  reg [15:0] codewords_120; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_185;
  reg [15:0] codewords_121; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_186;
  reg [15:0] codewords_122; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_187;
  reg [15:0] codewords_123; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_188;
  reg [15:0] codewords_124; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_189;
  reg [15:0] codewords_125; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_190;
  reg [15:0] codewords_126; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_191;
  reg [15:0] codewords_127; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_192;
  reg [15:0] codewords_128; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_193;
  reg [15:0] codewords_129; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_194;
  reg [15:0] codewords_130; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_195;
  reg [15:0] codewords_131; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_196;
  reg [15:0] codewords_132; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_197;
  reg [15:0] codewords_133; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_198;
  reg [15:0] codewords_134; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_199;
  reg [15:0] codewords_135; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_200;
  reg [15:0] codewords_136; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_201;
  reg [15:0] codewords_137; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_202;
  reg [15:0] codewords_138; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_203;
  reg [15:0] codewords_139; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_204;
  reg [15:0] codewords_140; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_205;
  reg [15:0] codewords_141; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_206;
  reg [15:0] codewords_142; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_207;
  reg [15:0] codewords_143; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_208;
  reg [15:0] codewords_144; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_209;
  reg [15:0] codewords_145; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_210;
  reg [15:0] codewords_146; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_211;
  reg [15:0] codewords_147; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_212;
  reg [15:0] codewords_148; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_213;
  reg [15:0] codewords_149; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_214;
  reg [15:0] codewords_150; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_215;
  reg [15:0] codewords_151; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_216;
  reg [15:0] codewords_152; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_217;
  reg [15:0] codewords_153; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_218;
  reg [15:0] codewords_154; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_219;
  reg [15:0] codewords_155; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_220;
  reg [15:0] codewords_156; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_221;
  reg [15:0] codewords_157; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_222;
  reg [15:0] codewords_158; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_223;
  reg [15:0] codewords_159; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_224;
  reg [15:0] codewords_160; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_225;
  reg [15:0] codewords_161; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_226;
  reg [15:0] codewords_162; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_227;
  reg [15:0] codewords_163; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_228;
  reg [15:0] codewords_164; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_229;
  reg [15:0] codewords_165; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_230;
  reg [15:0] codewords_166; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_231;
  reg [15:0] codewords_167; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_232;
  reg [15:0] codewords_168; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_233;
  reg [15:0] codewords_169; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_234;
  reg [15:0] codewords_170; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_235;
  reg [15:0] codewords_171; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_236;
  reg [15:0] codewords_172; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_237;
  reg [15:0] codewords_173; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_238;
  reg [15:0] codewords_174; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_239;
  reg [15:0] codewords_175; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_240;
  reg [15:0] codewords_176; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_241;
  reg [15:0] codewords_177; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_242;
  reg [15:0] codewords_178; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_243;
  reg [15:0] codewords_179; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_244;
  reg [15:0] codewords_180; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_245;
  reg [15:0] codewords_181; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_246;
  reg [15:0] codewords_182; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_247;
  reg [15:0] codewords_183; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_248;
  reg [15:0] codewords_184; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_249;
  reg [15:0] codewords_185; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_250;
  reg [15:0] codewords_186; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_251;
  reg [15:0] codewords_187; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_252;
  reg [15:0] codewords_188; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_253;
  reg [15:0] codewords_189; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_254;
  reg [15:0] codewords_190; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_255;
  reg [15:0] codewords_191; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_256;
  reg [15:0] codewords_192; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_257;
  reg [15:0] codewords_193; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_258;
  reg [15:0] codewords_194; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_259;
  reg [15:0] codewords_195; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_260;
  reg [15:0] codewords_196; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_261;
  reg [15:0] codewords_197; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_262;
  reg [15:0] codewords_198; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_263;
  reg [15:0] codewords_199; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_264;
  reg [15:0] codewords_200; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_265;
  reg [15:0] codewords_201; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_266;
  reg [15:0] codewords_202; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_267;
  reg [15:0] codewords_203; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_268;
  reg [15:0] codewords_204; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_269;
  reg [15:0] codewords_205; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_270;
  reg [15:0] codewords_206; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_271;
  reg [15:0] codewords_207; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_272;
  reg [15:0] codewords_208; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_273;
  reg [15:0] codewords_209; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_274;
  reg [15:0] codewords_210; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_275;
  reg [15:0] codewords_211; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_276;
  reg [15:0] codewords_212; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_277;
  reg [15:0] codewords_213; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_278;
  reg [15:0] codewords_214; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_279;
  reg [15:0] codewords_215; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_280;
  reg [15:0] codewords_216; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_281;
  reg [15:0] codewords_217; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_282;
  reg [15:0] codewords_218; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_283;
  reg [15:0] codewords_219; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_284;
  reg [15:0] codewords_220; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_285;
  reg [15:0] codewords_221; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_286;
  reg [15:0] codewords_222; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_287;
  reg [15:0] codewords_223; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_288;
  reg [15:0] codewords_224; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_289;
  reg [15:0] codewords_225; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_290;
  reg [15:0] codewords_226; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_291;
  reg [15:0] codewords_227; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_292;
  reg [15:0] codewords_228; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_293;
  reg [15:0] codewords_229; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_294;
  reg [15:0] codewords_230; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_295;
  reg [15:0] codewords_231; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_296;
  reg [15:0] codewords_232; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_297;
  reg [15:0] codewords_233; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_298;
  reg [15:0] codewords_234; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_299;
  reg [15:0] codewords_235; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_300;
  reg [15:0] codewords_236; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_301;
  reg [15:0] codewords_237; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_302;
  reg [15:0] codewords_238; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_303;
  reg [15:0] codewords_239; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_304;
  reg [15:0] codewords_240; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_305;
  reg [15:0] codewords_241; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_306;
  reg [15:0] codewords_242; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_307;
  reg [15:0] codewords_243; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_308;
  reg [15:0] codewords_244; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_309;
  reg [15:0] codewords_245; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_310;
  reg [15:0] codewords_246; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_311;
  reg [15:0] codewords_247; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_312;
  reg [15:0] codewords_248; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_313;
  reg [15:0] codewords_249; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_314;
  reg [15:0] codewords_250; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_315;
  reg [15:0] codewords_251; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_316;
  reg [15:0] codewords_252; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_317;
  reg [15:0] codewords_253; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_318;
  reg [15:0] codewords_254; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_319;
  reg [15:0] codewords_255; // @[codewordGenerator.scala 46:26]
  reg [31:0] _RAND_320;
  reg [23:0] codewordsOut_0; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_321;
  reg [23:0] codewordsOut_1; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_322;
  reg [23:0] codewordsOut_2; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_323;
  reg [23:0] codewordsOut_3; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_324;
  reg [23:0] codewordsOut_4; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_325;
  reg [23:0] codewordsOut_5; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_326;
  reg [23:0] codewordsOut_6; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_327;
  reg [23:0] codewordsOut_7; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_328;
  reg [23:0] codewordsOut_8; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_329;
  reg [23:0] codewordsOut_9; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_330;
  reg [23:0] codewordsOut_10; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_331;
  reg [23:0] codewordsOut_11; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_332;
  reg [23:0] codewordsOut_12; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_333;
  reg [23:0] codewordsOut_13; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_334;
  reg [23:0] codewordsOut_14; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_335;
  reg [23:0] codewordsOut_15; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_336;
  reg [23:0] codewordsOut_16; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_337;
  reg [23:0] codewordsOut_17; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_338;
  reg [23:0] codewordsOut_18; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_339;
  reg [23:0] codewordsOut_19; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_340;
  reg [23:0] codewordsOut_20; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_341;
  reg [23:0] codewordsOut_21; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_342;
  reg [23:0] codewordsOut_22; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_343;
  reg [23:0] codewordsOut_23; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_344;
  reg [23:0] codewordsOut_24; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_345;
  reg [23:0] codewordsOut_25; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_346;
  reg [23:0] codewordsOut_26; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_347;
  reg [23:0] codewordsOut_27; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_348;
  reg [23:0] codewordsOut_28; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_349;
  reg [23:0] codewordsOut_29; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_350;
  reg [23:0] codewordsOut_30; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_351;
  reg [23:0] codewordsOut_31; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_352;
  reg [23:0] codewordsOut_32; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_353;
  reg [23:0] codewordsOut_33; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_354;
  reg [23:0] codewordsOut_34; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_355;
  reg [23:0] codewordsOut_35; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_356;
  reg [23:0] codewordsOut_36; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_357;
  reg [23:0] codewordsOut_37; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_358;
  reg [23:0] codewordsOut_38; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_359;
  reg [23:0] codewordsOut_39; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_360;
  reg [23:0] codewordsOut_40; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_361;
  reg [23:0] codewordsOut_41; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_362;
  reg [23:0] codewordsOut_42; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_363;
  reg [23:0] codewordsOut_43; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_364;
  reg [23:0] codewordsOut_44; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_365;
  reg [23:0] codewordsOut_45; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_366;
  reg [23:0] codewordsOut_46; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_367;
  reg [23:0] codewordsOut_47; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_368;
  reg [23:0] codewordsOut_48; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_369;
  reg [23:0] codewordsOut_49; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_370;
  reg [23:0] codewordsOut_50; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_371;
  reg [23:0] codewordsOut_51; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_372;
  reg [23:0] codewordsOut_52; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_373;
  reg [23:0] codewordsOut_53; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_374;
  reg [23:0] codewordsOut_54; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_375;
  reg [23:0] codewordsOut_55; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_376;
  reg [23:0] codewordsOut_56; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_377;
  reg [23:0] codewordsOut_57; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_378;
  reg [23:0] codewordsOut_58; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_379;
  reg [23:0] codewordsOut_59; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_380;
  reg [23:0] codewordsOut_60; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_381;
  reg [23:0] codewordsOut_61; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_382;
  reg [23:0] codewordsOut_62; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_383;
  reg [23:0] codewordsOut_63; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_384;
  reg [23:0] codewordsOut_64; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_385;
  reg [23:0] codewordsOut_65; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_386;
  reg [23:0] codewordsOut_66; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_387;
  reg [23:0] codewordsOut_67; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_388;
  reg [23:0] codewordsOut_68; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_389;
  reg [23:0] codewordsOut_69; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_390;
  reg [23:0] codewordsOut_70; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_391;
  reg [23:0] codewordsOut_71; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_392;
  reg [23:0] codewordsOut_72; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_393;
  reg [23:0] codewordsOut_73; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_394;
  reg [23:0] codewordsOut_74; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_395;
  reg [23:0] codewordsOut_75; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_396;
  reg [23:0] codewordsOut_76; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_397;
  reg [23:0] codewordsOut_77; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_398;
  reg [23:0] codewordsOut_78; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_399;
  reg [23:0] codewordsOut_79; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_400;
  reg [23:0] codewordsOut_80; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_401;
  reg [23:0] codewordsOut_81; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_402;
  reg [23:0] codewordsOut_82; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_403;
  reg [23:0] codewordsOut_83; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_404;
  reg [23:0] codewordsOut_84; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_405;
  reg [23:0] codewordsOut_85; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_406;
  reg [23:0] codewordsOut_86; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_407;
  reg [23:0] codewordsOut_87; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_408;
  reg [23:0] codewordsOut_88; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_409;
  reg [23:0] codewordsOut_89; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_410;
  reg [23:0] codewordsOut_90; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_411;
  reg [23:0] codewordsOut_91; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_412;
  reg [23:0] codewordsOut_92; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_413;
  reg [23:0] codewordsOut_93; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_414;
  reg [23:0] codewordsOut_94; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_415;
  reg [23:0] codewordsOut_95; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_416;
  reg [23:0] codewordsOut_96; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_417;
  reg [23:0] codewordsOut_97; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_418;
  reg [23:0] codewordsOut_98; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_419;
  reg [23:0] codewordsOut_99; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_420;
  reg [23:0] codewordsOut_100; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_421;
  reg [23:0] codewordsOut_101; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_422;
  reg [23:0] codewordsOut_102; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_423;
  reg [23:0] codewordsOut_103; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_424;
  reg [23:0] codewordsOut_104; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_425;
  reg [23:0] codewordsOut_105; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_426;
  reg [23:0] codewordsOut_106; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_427;
  reg [23:0] codewordsOut_107; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_428;
  reg [23:0] codewordsOut_108; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_429;
  reg [23:0] codewordsOut_109; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_430;
  reg [23:0] codewordsOut_110; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_431;
  reg [23:0] codewordsOut_111; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_432;
  reg [23:0] codewordsOut_112; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_433;
  reg [23:0] codewordsOut_113; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_434;
  reg [23:0] codewordsOut_114; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_435;
  reg [23:0] codewordsOut_115; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_436;
  reg [23:0] codewordsOut_116; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_437;
  reg [23:0] codewordsOut_117; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_438;
  reg [23:0] codewordsOut_118; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_439;
  reg [23:0] codewordsOut_119; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_440;
  reg [23:0] codewordsOut_120; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_441;
  reg [23:0] codewordsOut_121; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_442;
  reg [23:0] codewordsOut_122; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_443;
  reg [23:0] codewordsOut_123; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_444;
  reg [23:0] codewordsOut_124; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_445;
  reg [23:0] codewordsOut_125; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_446;
  reg [23:0] codewordsOut_126; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_447;
  reg [23:0] codewordsOut_127; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_448;
  reg [23:0] codewordsOut_128; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_449;
  reg [23:0] codewordsOut_129; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_450;
  reg [23:0] codewordsOut_130; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_451;
  reg [23:0] codewordsOut_131; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_452;
  reg [23:0] codewordsOut_132; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_453;
  reg [23:0] codewordsOut_133; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_454;
  reg [23:0] codewordsOut_134; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_455;
  reg [23:0] codewordsOut_135; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_456;
  reg [23:0] codewordsOut_136; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_457;
  reg [23:0] codewordsOut_137; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_458;
  reg [23:0] codewordsOut_138; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_459;
  reg [23:0] codewordsOut_139; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_460;
  reg [23:0] codewordsOut_140; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_461;
  reg [23:0] codewordsOut_141; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_462;
  reg [23:0] codewordsOut_142; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_463;
  reg [23:0] codewordsOut_143; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_464;
  reg [23:0] codewordsOut_144; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_465;
  reg [23:0] codewordsOut_145; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_466;
  reg [23:0] codewordsOut_146; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_467;
  reg [23:0] codewordsOut_147; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_468;
  reg [23:0] codewordsOut_148; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_469;
  reg [23:0] codewordsOut_149; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_470;
  reg [23:0] codewordsOut_150; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_471;
  reg [23:0] codewordsOut_151; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_472;
  reg [23:0] codewordsOut_152; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_473;
  reg [23:0] codewordsOut_153; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_474;
  reg [23:0] codewordsOut_154; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_475;
  reg [23:0] codewordsOut_155; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_476;
  reg [23:0] codewordsOut_156; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_477;
  reg [23:0] codewordsOut_157; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_478;
  reg [23:0] codewordsOut_158; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_479;
  reg [23:0] codewordsOut_159; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_480;
  reg [23:0] codewordsOut_160; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_481;
  reg [23:0] codewordsOut_161; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_482;
  reg [23:0] codewordsOut_162; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_483;
  reg [23:0] codewordsOut_163; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_484;
  reg [23:0] codewordsOut_164; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_485;
  reg [23:0] codewordsOut_165; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_486;
  reg [23:0] codewordsOut_166; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_487;
  reg [23:0] codewordsOut_167; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_488;
  reg [23:0] codewordsOut_168; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_489;
  reg [23:0] codewordsOut_169; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_490;
  reg [23:0] codewordsOut_170; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_491;
  reg [23:0] codewordsOut_171; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_492;
  reg [23:0] codewordsOut_172; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_493;
  reg [23:0] codewordsOut_173; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_494;
  reg [23:0] codewordsOut_174; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_495;
  reg [23:0] codewordsOut_175; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_496;
  reg [23:0] codewordsOut_176; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_497;
  reg [23:0] codewordsOut_177; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_498;
  reg [23:0] codewordsOut_178; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_499;
  reg [23:0] codewordsOut_179; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_500;
  reg [23:0] codewordsOut_180; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_501;
  reg [23:0] codewordsOut_181; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_502;
  reg [23:0] codewordsOut_182; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_503;
  reg [23:0] codewordsOut_183; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_504;
  reg [23:0] codewordsOut_184; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_505;
  reg [23:0] codewordsOut_185; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_506;
  reg [23:0] codewordsOut_186; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_507;
  reg [23:0] codewordsOut_187; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_508;
  reg [23:0] codewordsOut_188; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_509;
  reg [23:0] codewordsOut_189; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_510;
  reg [23:0] codewordsOut_190; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_511;
  reg [23:0] codewordsOut_191; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_512;
  reg [23:0] codewordsOut_192; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_513;
  reg [23:0] codewordsOut_193; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_514;
  reg [23:0] codewordsOut_194; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_515;
  reg [23:0] codewordsOut_195; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_516;
  reg [23:0] codewordsOut_196; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_517;
  reg [23:0] codewordsOut_197; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_518;
  reg [23:0] codewordsOut_198; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_519;
  reg [23:0] codewordsOut_199; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_520;
  reg [23:0] codewordsOut_200; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_521;
  reg [23:0] codewordsOut_201; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_522;
  reg [23:0] codewordsOut_202; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_523;
  reg [23:0] codewordsOut_203; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_524;
  reg [23:0] codewordsOut_204; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_525;
  reg [23:0] codewordsOut_205; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_526;
  reg [23:0] codewordsOut_206; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_527;
  reg [23:0] codewordsOut_207; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_528;
  reg [23:0] codewordsOut_208; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_529;
  reg [23:0] codewordsOut_209; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_530;
  reg [23:0] codewordsOut_210; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_531;
  reg [23:0] codewordsOut_211; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_532;
  reg [23:0] codewordsOut_212; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_533;
  reg [23:0] codewordsOut_213; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_534;
  reg [23:0] codewordsOut_214; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_535;
  reg [23:0] codewordsOut_215; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_536;
  reg [23:0] codewordsOut_216; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_537;
  reg [23:0] codewordsOut_217; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_538;
  reg [23:0] codewordsOut_218; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_539;
  reg [23:0] codewordsOut_219; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_540;
  reg [23:0] codewordsOut_220; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_541;
  reg [23:0] codewordsOut_221; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_542;
  reg [23:0] codewordsOut_222; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_543;
  reg [23:0] codewordsOut_223; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_544;
  reg [23:0] codewordsOut_224; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_545;
  reg [23:0] codewordsOut_225; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_546;
  reg [23:0] codewordsOut_226; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_547;
  reg [23:0] codewordsOut_227; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_548;
  reg [23:0] codewordsOut_228; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_549;
  reg [23:0] codewordsOut_229; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_550;
  reg [23:0] codewordsOut_230; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_551;
  reg [23:0] codewordsOut_231; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_552;
  reg [23:0] codewordsOut_232; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_553;
  reg [23:0] codewordsOut_233; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_554;
  reg [23:0] codewordsOut_234; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_555;
  reg [23:0] codewordsOut_235; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_556;
  reg [23:0] codewordsOut_236; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_557;
  reg [23:0] codewordsOut_237; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_558;
  reg [23:0] codewordsOut_238; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_559;
  reg [23:0] codewordsOut_239; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_560;
  reg [23:0] codewordsOut_240; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_561;
  reg [23:0] codewordsOut_241; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_562;
  reg [23:0] codewordsOut_242; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_563;
  reg [23:0] codewordsOut_243; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_564;
  reg [23:0] codewordsOut_244; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_565;
  reg [23:0] codewordsOut_245; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_566;
  reg [23:0] codewordsOut_246; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_567;
  reg [23:0] codewordsOut_247; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_568;
  reg [23:0] codewordsOut_248; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_569;
  reg [23:0] codewordsOut_249; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_570;
  reg [23:0] codewordsOut_250; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_571;
  reg [23:0] codewordsOut_251; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_572;
  reg [23:0] codewordsOut_252; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_573;
  reg [23:0] codewordsOut_253; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_574;
  reg [23:0] codewordsOut_254; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_575;
  reg [23:0] codewordsOut_255; // @[codewordGenerator.scala 47:25]
  reg [31:0] _RAND_576;
  reg [4:0] lengths_0; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_577;
  reg [4:0] lengths_1; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_578;
  reg [4:0] lengths_2; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_579;
  reg [4:0] lengths_3; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_580;
  reg [4:0] lengths_4; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_581;
  reg [4:0] lengths_5; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_582;
  reg [4:0] lengths_6; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_583;
  reg [4:0] lengths_7; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_584;
  reg [4:0] lengths_8; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_585;
  reg [4:0] lengths_9; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_586;
  reg [4:0] lengths_10; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_587;
  reg [4:0] lengths_11; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_588;
  reg [4:0] lengths_12; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_589;
  reg [4:0] lengths_13; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_590;
  reg [4:0] lengths_14; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_591;
  reg [4:0] lengths_15; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_592;
  reg [4:0] lengths_16; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_593;
  reg [4:0] lengths_17; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_594;
  reg [4:0] lengths_18; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_595;
  reg [4:0] lengths_19; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_596;
  reg [4:0] lengths_20; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_597;
  reg [4:0] lengths_21; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_598;
  reg [4:0] lengths_22; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_599;
  reg [4:0] lengths_23; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_600;
  reg [4:0] lengths_24; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_601;
  reg [4:0] lengths_25; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_602;
  reg [4:0] lengths_26; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_603;
  reg [4:0] lengths_27; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_604;
  reg [4:0] lengths_28; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_605;
  reg [4:0] lengths_29; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_606;
  reg [4:0] lengths_30; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_607;
  reg [4:0] lengths_31; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_608;
  reg [4:0] lengths_32; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_609;
  reg [4:0] lengths_33; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_610;
  reg [4:0] lengths_34; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_611;
  reg [4:0] lengths_35; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_612;
  reg [4:0] lengths_36; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_613;
  reg [4:0] lengths_37; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_614;
  reg [4:0] lengths_38; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_615;
  reg [4:0] lengths_39; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_616;
  reg [4:0] lengths_40; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_617;
  reg [4:0] lengths_41; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_618;
  reg [4:0] lengths_42; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_619;
  reg [4:0] lengths_43; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_620;
  reg [4:0] lengths_44; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_621;
  reg [4:0] lengths_45; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_622;
  reg [4:0] lengths_46; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_623;
  reg [4:0] lengths_47; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_624;
  reg [4:0] lengths_48; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_625;
  reg [4:0] lengths_49; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_626;
  reg [4:0] lengths_50; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_627;
  reg [4:0] lengths_51; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_628;
  reg [4:0] lengths_52; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_629;
  reg [4:0] lengths_53; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_630;
  reg [4:0] lengths_54; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_631;
  reg [4:0] lengths_55; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_632;
  reg [4:0] lengths_56; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_633;
  reg [4:0] lengths_57; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_634;
  reg [4:0] lengths_58; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_635;
  reg [4:0] lengths_59; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_636;
  reg [4:0] lengths_60; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_637;
  reg [4:0] lengths_61; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_638;
  reg [4:0] lengths_62; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_639;
  reg [4:0] lengths_63; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_640;
  reg [4:0] lengths_64; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_641;
  reg [4:0] lengths_65; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_642;
  reg [4:0] lengths_66; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_643;
  reg [4:0] lengths_67; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_644;
  reg [4:0] lengths_68; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_645;
  reg [4:0] lengths_69; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_646;
  reg [4:0] lengths_70; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_647;
  reg [4:0] lengths_71; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_648;
  reg [4:0] lengths_72; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_649;
  reg [4:0] lengths_73; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_650;
  reg [4:0] lengths_74; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_651;
  reg [4:0] lengths_75; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_652;
  reg [4:0] lengths_76; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_653;
  reg [4:0] lengths_77; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_654;
  reg [4:0] lengths_78; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_655;
  reg [4:0] lengths_79; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_656;
  reg [4:0] lengths_80; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_657;
  reg [4:0] lengths_81; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_658;
  reg [4:0] lengths_82; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_659;
  reg [4:0] lengths_83; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_660;
  reg [4:0] lengths_84; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_661;
  reg [4:0] lengths_85; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_662;
  reg [4:0] lengths_86; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_663;
  reg [4:0] lengths_87; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_664;
  reg [4:0] lengths_88; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_665;
  reg [4:0] lengths_89; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_666;
  reg [4:0] lengths_90; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_667;
  reg [4:0] lengths_91; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_668;
  reg [4:0] lengths_92; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_669;
  reg [4:0] lengths_93; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_670;
  reg [4:0] lengths_94; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_671;
  reg [4:0] lengths_95; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_672;
  reg [4:0] lengths_96; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_673;
  reg [4:0] lengths_97; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_674;
  reg [4:0] lengths_98; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_675;
  reg [4:0] lengths_99; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_676;
  reg [4:0] lengths_100; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_677;
  reg [4:0] lengths_101; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_678;
  reg [4:0] lengths_102; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_679;
  reg [4:0] lengths_103; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_680;
  reg [4:0] lengths_104; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_681;
  reg [4:0] lengths_105; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_682;
  reg [4:0] lengths_106; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_683;
  reg [4:0] lengths_107; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_684;
  reg [4:0] lengths_108; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_685;
  reg [4:0] lengths_109; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_686;
  reg [4:0] lengths_110; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_687;
  reg [4:0] lengths_111; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_688;
  reg [4:0] lengths_112; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_689;
  reg [4:0] lengths_113; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_690;
  reg [4:0] lengths_114; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_691;
  reg [4:0] lengths_115; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_692;
  reg [4:0] lengths_116; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_693;
  reg [4:0] lengths_117; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_694;
  reg [4:0] lengths_118; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_695;
  reg [4:0] lengths_119; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_696;
  reg [4:0] lengths_120; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_697;
  reg [4:0] lengths_121; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_698;
  reg [4:0] lengths_122; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_699;
  reg [4:0] lengths_123; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_700;
  reg [4:0] lengths_124; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_701;
  reg [4:0] lengths_125; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_702;
  reg [4:0] lengths_126; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_703;
  reg [4:0] lengths_127; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_704;
  reg [4:0] lengths_128; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_705;
  reg [4:0] lengths_129; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_706;
  reg [4:0] lengths_130; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_707;
  reg [4:0] lengths_131; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_708;
  reg [4:0] lengths_132; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_709;
  reg [4:0] lengths_133; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_710;
  reg [4:0] lengths_134; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_711;
  reg [4:0] lengths_135; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_712;
  reg [4:0] lengths_136; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_713;
  reg [4:0] lengths_137; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_714;
  reg [4:0] lengths_138; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_715;
  reg [4:0] lengths_139; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_716;
  reg [4:0] lengths_140; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_717;
  reg [4:0] lengths_141; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_718;
  reg [4:0] lengths_142; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_719;
  reg [4:0] lengths_143; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_720;
  reg [4:0] lengths_144; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_721;
  reg [4:0] lengths_145; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_722;
  reg [4:0] lengths_146; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_723;
  reg [4:0] lengths_147; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_724;
  reg [4:0] lengths_148; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_725;
  reg [4:0] lengths_149; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_726;
  reg [4:0] lengths_150; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_727;
  reg [4:0] lengths_151; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_728;
  reg [4:0] lengths_152; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_729;
  reg [4:0] lengths_153; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_730;
  reg [4:0] lengths_154; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_731;
  reg [4:0] lengths_155; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_732;
  reg [4:0] lengths_156; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_733;
  reg [4:0] lengths_157; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_734;
  reg [4:0] lengths_158; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_735;
  reg [4:0] lengths_159; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_736;
  reg [4:0] lengths_160; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_737;
  reg [4:0] lengths_161; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_738;
  reg [4:0] lengths_162; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_739;
  reg [4:0] lengths_163; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_740;
  reg [4:0] lengths_164; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_741;
  reg [4:0] lengths_165; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_742;
  reg [4:0] lengths_166; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_743;
  reg [4:0] lengths_167; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_744;
  reg [4:0] lengths_168; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_745;
  reg [4:0] lengths_169; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_746;
  reg [4:0] lengths_170; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_747;
  reg [4:0] lengths_171; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_748;
  reg [4:0] lengths_172; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_749;
  reg [4:0] lengths_173; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_750;
  reg [4:0] lengths_174; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_751;
  reg [4:0] lengths_175; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_752;
  reg [4:0] lengths_176; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_753;
  reg [4:0] lengths_177; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_754;
  reg [4:0] lengths_178; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_755;
  reg [4:0] lengths_179; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_756;
  reg [4:0] lengths_180; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_757;
  reg [4:0] lengths_181; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_758;
  reg [4:0] lengths_182; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_759;
  reg [4:0] lengths_183; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_760;
  reg [4:0] lengths_184; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_761;
  reg [4:0] lengths_185; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_762;
  reg [4:0] lengths_186; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_763;
  reg [4:0] lengths_187; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_764;
  reg [4:0] lengths_188; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_765;
  reg [4:0] lengths_189; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_766;
  reg [4:0] lengths_190; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_767;
  reg [4:0] lengths_191; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_768;
  reg [4:0] lengths_192; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_769;
  reg [4:0] lengths_193; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_770;
  reg [4:0] lengths_194; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_771;
  reg [4:0] lengths_195; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_772;
  reg [4:0] lengths_196; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_773;
  reg [4:0] lengths_197; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_774;
  reg [4:0] lengths_198; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_775;
  reg [4:0] lengths_199; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_776;
  reg [4:0] lengths_200; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_777;
  reg [4:0] lengths_201; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_778;
  reg [4:0] lengths_202; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_779;
  reg [4:0] lengths_203; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_780;
  reg [4:0] lengths_204; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_781;
  reg [4:0] lengths_205; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_782;
  reg [4:0] lengths_206; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_783;
  reg [4:0] lengths_207; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_784;
  reg [4:0] lengths_208; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_785;
  reg [4:0] lengths_209; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_786;
  reg [4:0] lengths_210; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_787;
  reg [4:0] lengths_211; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_788;
  reg [4:0] lengths_212; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_789;
  reg [4:0] lengths_213; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_790;
  reg [4:0] lengths_214; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_791;
  reg [4:0] lengths_215; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_792;
  reg [4:0] lengths_216; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_793;
  reg [4:0] lengths_217; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_794;
  reg [4:0] lengths_218; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_795;
  reg [4:0] lengths_219; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_796;
  reg [4:0] lengths_220; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_797;
  reg [4:0] lengths_221; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_798;
  reg [4:0] lengths_222; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_799;
  reg [4:0] lengths_223; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_800;
  reg [4:0] lengths_224; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_801;
  reg [4:0] lengths_225; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_802;
  reg [4:0] lengths_226; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_803;
  reg [4:0] lengths_227; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_804;
  reg [4:0] lengths_228; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_805;
  reg [4:0] lengths_229; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_806;
  reg [4:0] lengths_230; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_807;
  reg [4:0] lengths_231; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_808;
  reg [4:0] lengths_232; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_809;
  reg [4:0] lengths_233; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_810;
  reg [4:0] lengths_234; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_811;
  reg [4:0] lengths_235; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_812;
  reg [4:0] lengths_236; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_813;
  reg [4:0] lengths_237; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_814;
  reg [4:0] lengths_238; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_815;
  reg [4:0] lengths_239; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_816;
  reg [4:0] lengths_240; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_817;
  reg [4:0] lengths_241; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_818;
  reg [4:0] lengths_242; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_819;
  reg [4:0] lengths_243; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_820;
  reg [4:0] lengths_244; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_821;
  reg [4:0] lengths_245; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_822;
  reg [4:0] lengths_246; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_823;
  reg [4:0] lengths_247; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_824;
  reg [4:0] lengths_248; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_825;
  reg [4:0] lengths_249; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_826;
  reg [4:0] lengths_250; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_827;
  reg [4:0] lengths_251; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_828;
  reg [4:0] lengths_252; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_829;
  reg [4:0] lengths_253; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_830;
  reg [4:0] lengths_254; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_831;
  reg [4:0] lengths_255; // @[codewordGenerator.scala 48:24]
  reg [31:0] _RAND_832;
  reg [4:0] lengthsOut_0; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_833;
  reg [4:0] lengthsOut_1; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_834;
  reg [4:0] lengthsOut_2; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_835;
  reg [4:0] lengthsOut_3; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_836;
  reg [4:0] lengthsOut_4; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_837;
  reg [4:0] lengthsOut_5; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_838;
  reg [4:0] lengthsOut_6; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_839;
  reg [4:0] lengthsOut_7; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_840;
  reg [4:0] lengthsOut_8; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_841;
  reg [4:0] lengthsOut_9; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_842;
  reg [4:0] lengthsOut_10; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_843;
  reg [4:0] lengthsOut_11; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_844;
  reg [4:0] lengthsOut_12; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_845;
  reg [4:0] lengthsOut_13; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_846;
  reg [4:0] lengthsOut_14; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_847;
  reg [4:0] lengthsOut_15; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_848;
  reg [4:0] lengthsOut_16; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_849;
  reg [4:0] lengthsOut_17; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_850;
  reg [4:0] lengthsOut_18; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_851;
  reg [4:0] lengthsOut_19; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_852;
  reg [4:0] lengthsOut_20; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_853;
  reg [4:0] lengthsOut_21; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_854;
  reg [4:0] lengthsOut_22; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_855;
  reg [4:0] lengthsOut_23; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_856;
  reg [4:0] lengthsOut_24; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_857;
  reg [4:0] lengthsOut_25; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_858;
  reg [4:0] lengthsOut_26; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_859;
  reg [4:0] lengthsOut_27; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_860;
  reg [4:0] lengthsOut_28; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_861;
  reg [4:0] lengthsOut_29; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_862;
  reg [4:0] lengthsOut_30; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_863;
  reg [4:0] lengthsOut_31; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_864;
  reg [4:0] lengthsOut_32; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_865;
  reg [4:0] lengthsOut_33; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_866;
  reg [4:0] lengthsOut_34; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_867;
  reg [4:0] lengthsOut_35; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_868;
  reg [4:0] lengthsOut_36; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_869;
  reg [4:0] lengthsOut_37; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_870;
  reg [4:0] lengthsOut_38; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_871;
  reg [4:0] lengthsOut_39; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_872;
  reg [4:0] lengthsOut_40; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_873;
  reg [4:0] lengthsOut_41; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_874;
  reg [4:0] lengthsOut_42; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_875;
  reg [4:0] lengthsOut_43; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_876;
  reg [4:0] lengthsOut_44; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_877;
  reg [4:0] lengthsOut_45; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_878;
  reg [4:0] lengthsOut_46; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_879;
  reg [4:0] lengthsOut_47; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_880;
  reg [4:0] lengthsOut_48; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_881;
  reg [4:0] lengthsOut_49; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_882;
  reg [4:0] lengthsOut_50; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_883;
  reg [4:0] lengthsOut_51; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_884;
  reg [4:0] lengthsOut_52; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_885;
  reg [4:0] lengthsOut_53; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_886;
  reg [4:0] lengthsOut_54; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_887;
  reg [4:0] lengthsOut_55; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_888;
  reg [4:0] lengthsOut_56; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_889;
  reg [4:0] lengthsOut_57; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_890;
  reg [4:0] lengthsOut_58; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_891;
  reg [4:0] lengthsOut_59; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_892;
  reg [4:0] lengthsOut_60; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_893;
  reg [4:0] lengthsOut_61; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_894;
  reg [4:0] lengthsOut_62; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_895;
  reg [4:0] lengthsOut_63; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_896;
  reg [4:0] lengthsOut_64; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_897;
  reg [4:0] lengthsOut_65; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_898;
  reg [4:0] lengthsOut_66; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_899;
  reg [4:0] lengthsOut_67; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_900;
  reg [4:0] lengthsOut_68; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_901;
  reg [4:0] lengthsOut_69; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_902;
  reg [4:0] lengthsOut_70; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_903;
  reg [4:0] lengthsOut_71; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_904;
  reg [4:0] lengthsOut_72; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_905;
  reg [4:0] lengthsOut_73; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_906;
  reg [4:0] lengthsOut_74; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_907;
  reg [4:0] lengthsOut_75; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_908;
  reg [4:0] lengthsOut_76; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_909;
  reg [4:0] lengthsOut_77; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_910;
  reg [4:0] lengthsOut_78; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_911;
  reg [4:0] lengthsOut_79; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_912;
  reg [4:0] lengthsOut_80; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_913;
  reg [4:0] lengthsOut_81; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_914;
  reg [4:0] lengthsOut_82; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_915;
  reg [4:0] lengthsOut_83; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_916;
  reg [4:0] lengthsOut_84; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_917;
  reg [4:0] lengthsOut_85; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_918;
  reg [4:0] lengthsOut_86; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_919;
  reg [4:0] lengthsOut_87; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_920;
  reg [4:0] lengthsOut_88; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_921;
  reg [4:0] lengthsOut_89; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_922;
  reg [4:0] lengthsOut_90; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_923;
  reg [4:0] lengthsOut_91; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_924;
  reg [4:0] lengthsOut_92; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_925;
  reg [4:0] lengthsOut_93; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_926;
  reg [4:0] lengthsOut_94; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_927;
  reg [4:0] lengthsOut_95; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_928;
  reg [4:0] lengthsOut_96; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_929;
  reg [4:0] lengthsOut_97; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_930;
  reg [4:0] lengthsOut_98; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_931;
  reg [4:0] lengthsOut_99; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_932;
  reg [4:0] lengthsOut_100; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_933;
  reg [4:0] lengthsOut_101; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_934;
  reg [4:0] lengthsOut_102; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_935;
  reg [4:0] lengthsOut_103; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_936;
  reg [4:0] lengthsOut_104; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_937;
  reg [4:0] lengthsOut_105; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_938;
  reg [4:0] lengthsOut_106; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_939;
  reg [4:0] lengthsOut_107; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_940;
  reg [4:0] lengthsOut_108; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_941;
  reg [4:0] lengthsOut_109; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_942;
  reg [4:0] lengthsOut_110; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_943;
  reg [4:0] lengthsOut_111; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_944;
  reg [4:0] lengthsOut_112; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_945;
  reg [4:0] lengthsOut_113; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_946;
  reg [4:0] lengthsOut_114; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_947;
  reg [4:0] lengthsOut_115; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_948;
  reg [4:0] lengthsOut_116; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_949;
  reg [4:0] lengthsOut_117; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_950;
  reg [4:0] lengthsOut_118; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_951;
  reg [4:0] lengthsOut_119; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_952;
  reg [4:0] lengthsOut_120; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_953;
  reg [4:0] lengthsOut_121; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_954;
  reg [4:0] lengthsOut_122; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_955;
  reg [4:0] lengthsOut_123; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_956;
  reg [4:0] lengthsOut_124; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_957;
  reg [4:0] lengthsOut_125; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_958;
  reg [4:0] lengthsOut_126; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_959;
  reg [4:0] lengthsOut_127; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_960;
  reg [4:0] lengthsOut_128; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_961;
  reg [4:0] lengthsOut_129; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_962;
  reg [4:0] lengthsOut_130; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_963;
  reg [4:0] lengthsOut_131; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_964;
  reg [4:0] lengthsOut_132; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_965;
  reg [4:0] lengthsOut_133; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_966;
  reg [4:0] lengthsOut_134; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_967;
  reg [4:0] lengthsOut_135; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_968;
  reg [4:0] lengthsOut_136; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_969;
  reg [4:0] lengthsOut_137; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_970;
  reg [4:0] lengthsOut_138; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_971;
  reg [4:0] lengthsOut_139; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_972;
  reg [4:0] lengthsOut_140; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_973;
  reg [4:0] lengthsOut_141; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_974;
  reg [4:0] lengthsOut_142; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_975;
  reg [4:0] lengthsOut_143; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_976;
  reg [4:0] lengthsOut_144; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_977;
  reg [4:0] lengthsOut_145; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_978;
  reg [4:0] lengthsOut_146; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_979;
  reg [4:0] lengthsOut_147; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_980;
  reg [4:0] lengthsOut_148; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_981;
  reg [4:0] lengthsOut_149; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_982;
  reg [4:0] lengthsOut_150; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_983;
  reg [4:0] lengthsOut_151; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_984;
  reg [4:0] lengthsOut_152; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_985;
  reg [4:0] lengthsOut_153; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_986;
  reg [4:0] lengthsOut_154; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_987;
  reg [4:0] lengthsOut_155; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_988;
  reg [4:0] lengthsOut_156; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_989;
  reg [4:0] lengthsOut_157; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_990;
  reg [4:0] lengthsOut_158; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_991;
  reg [4:0] lengthsOut_159; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_992;
  reg [4:0] lengthsOut_160; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_993;
  reg [4:0] lengthsOut_161; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_994;
  reg [4:0] lengthsOut_162; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_995;
  reg [4:0] lengthsOut_163; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_996;
  reg [4:0] lengthsOut_164; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_997;
  reg [4:0] lengthsOut_165; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_998;
  reg [4:0] lengthsOut_166; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_999;
  reg [4:0] lengthsOut_167; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1000;
  reg [4:0] lengthsOut_168; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1001;
  reg [4:0] lengthsOut_169; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1002;
  reg [4:0] lengthsOut_170; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1003;
  reg [4:0] lengthsOut_171; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1004;
  reg [4:0] lengthsOut_172; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1005;
  reg [4:0] lengthsOut_173; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1006;
  reg [4:0] lengthsOut_174; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1007;
  reg [4:0] lengthsOut_175; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1008;
  reg [4:0] lengthsOut_176; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1009;
  reg [4:0] lengthsOut_177; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1010;
  reg [4:0] lengthsOut_178; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1011;
  reg [4:0] lengthsOut_179; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1012;
  reg [4:0] lengthsOut_180; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1013;
  reg [4:0] lengthsOut_181; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1014;
  reg [4:0] lengthsOut_182; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1015;
  reg [4:0] lengthsOut_183; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1016;
  reg [4:0] lengthsOut_184; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1017;
  reg [4:0] lengthsOut_185; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1018;
  reg [4:0] lengthsOut_186; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1019;
  reg [4:0] lengthsOut_187; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1020;
  reg [4:0] lengthsOut_188; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1021;
  reg [4:0] lengthsOut_189; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1022;
  reg [4:0] lengthsOut_190; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1023;
  reg [4:0] lengthsOut_191; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1024;
  reg [4:0] lengthsOut_192; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1025;
  reg [4:0] lengthsOut_193; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1026;
  reg [4:0] lengthsOut_194; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1027;
  reg [4:0] lengthsOut_195; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1028;
  reg [4:0] lengthsOut_196; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1029;
  reg [4:0] lengthsOut_197; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1030;
  reg [4:0] lengthsOut_198; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1031;
  reg [4:0] lengthsOut_199; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1032;
  reg [4:0] lengthsOut_200; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1033;
  reg [4:0] lengthsOut_201; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1034;
  reg [4:0] lengthsOut_202; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1035;
  reg [4:0] lengthsOut_203; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1036;
  reg [4:0] lengthsOut_204; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1037;
  reg [4:0] lengthsOut_205; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1038;
  reg [4:0] lengthsOut_206; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1039;
  reg [4:0] lengthsOut_207; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1040;
  reg [4:0] lengthsOut_208; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1041;
  reg [4:0] lengthsOut_209; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1042;
  reg [4:0] lengthsOut_210; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1043;
  reg [4:0] lengthsOut_211; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1044;
  reg [4:0] lengthsOut_212; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1045;
  reg [4:0] lengthsOut_213; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1046;
  reg [4:0] lengthsOut_214; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1047;
  reg [4:0] lengthsOut_215; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1048;
  reg [4:0] lengthsOut_216; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1049;
  reg [4:0] lengthsOut_217; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1050;
  reg [4:0] lengthsOut_218; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1051;
  reg [4:0] lengthsOut_219; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1052;
  reg [4:0] lengthsOut_220; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1053;
  reg [4:0] lengthsOut_221; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1054;
  reg [4:0] lengthsOut_222; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1055;
  reg [4:0] lengthsOut_223; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1056;
  reg [4:0] lengthsOut_224; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1057;
  reg [4:0] lengthsOut_225; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1058;
  reg [4:0] lengthsOut_226; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1059;
  reg [4:0] lengthsOut_227; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1060;
  reg [4:0] lengthsOut_228; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1061;
  reg [4:0] lengthsOut_229; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1062;
  reg [4:0] lengthsOut_230; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1063;
  reg [4:0] lengthsOut_231; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1064;
  reg [4:0] lengthsOut_232; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1065;
  reg [4:0] lengthsOut_233; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1066;
  reg [4:0] lengthsOut_234; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1067;
  reg [4:0] lengthsOut_235; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1068;
  reg [4:0] lengthsOut_236; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1069;
  reg [4:0] lengthsOut_237; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1070;
  reg [4:0] lengthsOut_238; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1071;
  reg [4:0] lengthsOut_239; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1072;
  reg [4:0] lengthsOut_240; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1073;
  reg [4:0] lengthsOut_241; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1074;
  reg [4:0] lengthsOut_242; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1075;
  reg [4:0] lengthsOut_243; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1076;
  reg [4:0] lengthsOut_244; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1077;
  reg [4:0] lengthsOut_245; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1078;
  reg [4:0] lengthsOut_246; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1079;
  reg [4:0] lengthsOut_247; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1080;
  reg [4:0] lengthsOut_248; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1081;
  reg [4:0] lengthsOut_249; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1082;
  reg [4:0] lengthsOut_250; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1083;
  reg [4:0] lengthsOut_251; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1084;
  reg [4:0] lengthsOut_252; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1085;
  reg [4:0] lengthsOut_253; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1086;
  reg [4:0] lengthsOut_254; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1087;
  reg [4:0] lengthsOut_255; // @[codewordGenerator.scala 49:23]
  reg [31:0] _RAND_1088;
  reg [7:0] characterIndex; // @[codewordGenerator.scala 51:31]
  reg [31:0] _RAND_1089;
  reg [8:0] nodes; // @[codewordGenerator.scala 52:22]
  reg [31:0] _RAND_1090;
  reg [3:0] characterDepth; // @[codewordGenerator.scala 53:31]
  reg [31:0] _RAND_1091;
  reg [15:0] codeword; // @[codewordGenerator.scala 54:25]
  reg [31:0] _RAND_1092;
  reg [15:0] escapeCodeword; // @[codewordGenerator.scala 55:31]
  reg [31:0] _RAND_1093;
  reg [3:0] escapeCharacterLength; // @[codewordGenerator.scala 57:38]
  reg [31:0] _RAND_1094;
  wire  _T_6 = state == 2'h0; // @[codewordGenerator.scala 63:14]
  wire [7:0] _GEN_33 = io_start ? io_inputs_depthsOut_0 : {{4'd0}, depths_0}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_34 = io_start ? io_inputs_depthsOut_1 : {{4'd0}, depths_1}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_35 = io_start ? io_inputs_depthsOut_2 : {{4'd0}, depths_2}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_36 = io_start ? io_inputs_depthsOut_3 : {{4'd0}, depths_3}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_37 = io_start ? io_inputs_depthsOut_4 : {{4'd0}, depths_4}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_38 = io_start ? io_inputs_depthsOut_5 : {{4'd0}, depths_5}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_39 = io_start ? io_inputs_depthsOut_6 : {{4'd0}, depths_6}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_40 = io_start ? io_inputs_depthsOut_7 : {{4'd0}, depths_7}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_41 = io_start ? io_inputs_depthsOut_8 : {{4'd0}, depths_8}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_42 = io_start ? io_inputs_depthsOut_9 : {{4'd0}, depths_9}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_43 = io_start ? io_inputs_depthsOut_10 : {{4'd0}, depths_10}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_44 = io_start ? io_inputs_depthsOut_11 : {{4'd0}, depths_11}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_45 = io_start ? io_inputs_depthsOut_12 : {{4'd0}, depths_12}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_46 = io_start ? io_inputs_depthsOut_13 : {{4'd0}, depths_13}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_47 = io_start ? io_inputs_depthsOut_14 : {{4'd0}, depths_14}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_48 = io_start ? io_inputs_depthsOut_15 : {{4'd0}, depths_15}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_49 = io_start ? io_inputs_depthsOut_16 : {{4'd0}, depths_16}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_50 = io_start ? io_inputs_depthsOut_17 : {{4'd0}, depths_17}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_51 = io_start ? io_inputs_depthsOut_18 : {{4'd0}, depths_18}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_52 = io_start ? io_inputs_depthsOut_19 : {{4'd0}, depths_19}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_53 = io_start ? io_inputs_depthsOut_20 : {{4'd0}, depths_20}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_54 = io_start ? io_inputs_depthsOut_21 : {{4'd0}, depths_21}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_55 = io_start ? io_inputs_depthsOut_22 : {{4'd0}, depths_22}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_56 = io_start ? io_inputs_depthsOut_23 : {{4'd0}, depths_23}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_57 = io_start ? io_inputs_depthsOut_24 : {{4'd0}, depths_24}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_58 = io_start ? io_inputs_depthsOut_25 : {{4'd0}, depths_25}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_59 = io_start ? io_inputs_depthsOut_26 : {{4'd0}, depths_26}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_60 = io_start ? io_inputs_depthsOut_27 : {{4'd0}, depths_27}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_61 = io_start ? io_inputs_depthsOut_28 : {{4'd0}, depths_28}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_62 = io_start ? io_inputs_depthsOut_29 : {{4'd0}, depths_29}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_63 = io_start ? io_inputs_depthsOut_30 : {{4'd0}, depths_30}; // @[codewordGenerator.scala 64:31]
  wire [7:0] _GEN_64 = io_start ? io_inputs_depthsOut_31 : {{4'd0}, depths_31}; // @[codewordGenerator.scala 64:31]
  wire [15:0] _GEN_84 = io_start ? 16'h0 : codeword; // @[codewordGenerator.scala 64:31]
  wire  _T_9 = state == 2'h1; // @[codewordGenerator.scala 76:20]
  wire [7:0] _T_12 = characterIndex + 8'h1; // @[codewordGenerator.scala 79:61]
  wire [3:0] _GEN_88 = 5'h1 == characterIndex[4:0] ? depths_1 : depths_0; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_89 = 5'h2 == characterIndex[4:0] ? depths_2 : _GEN_88; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_90 = 5'h3 == characterIndex[4:0] ? depths_3 : _GEN_89; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_91 = 5'h4 == characterIndex[4:0] ? depths_4 : _GEN_90; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_92 = 5'h5 == characterIndex[4:0] ? depths_5 : _GEN_91; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_93 = 5'h6 == characterIndex[4:0] ? depths_6 : _GEN_92; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_94 = 5'h7 == characterIndex[4:0] ? depths_7 : _GEN_93; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_95 = 5'h8 == characterIndex[4:0] ? depths_8 : _GEN_94; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_96 = 5'h9 == characterIndex[4:0] ? depths_9 : _GEN_95; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_97 = 5'ha == characterIndex[4:0] ? depths_10 : _GEN_96; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_98 = 5'hb == characterIndex[4:0] ? depths_11 : _GEN_97; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_99 = 5'hc == characterIndex[4:0] ? depths_12 : _GEN_98; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_100 = 5'hd == characterIndex[4:0] ? depths_13 : _GEN_99; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_101 = 5'he == characterIndex[4:0] ? depths_14 : _GEN_100; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_102 = 5'hf == characterIndex[4:0] ? depths_15 : _GEN_101; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_103 = 5'h10 == characterIndex[4:0] ? depths_16 : _GEN_102; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_104 = 5'h11 == characterIndex[4:0] ? depths_17 : _GEN_103; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_105 = 5'h12 == characterIndex[4:0] ? depths_18 : _GEN_104; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_106 = 5'h13 == characterIndex[4:0] ? depths_19 : _GEN_105; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_107 = 5'h14 == characterIndex[4:0] ? depths_20 : _GEN_106; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_108 = 5'h15 == characterIndex[4:0] ? depths_21 : _GEN_107; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_109 = 5'h16 == characterIndex[4:0] ? depths_22 : _GEN_108; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_110 = 5'h17 == characterIndex[4:0] ? depths_23 : _GEN_109; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_111 = 5'h18 == characterIndex[4:0] ? depths_24 : _GEN_110; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_112 = 5'h19 == characterIndex[4:0] ? depths_25 : _GEN_111; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_113 = 5'h1a == characterIndex[4:0] ? depths_26 : _GEN_112; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_114 = 5'h1b == characterIndex[4:0] ? depths_27 : _GEN_113; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_115 = 5'h1c == characterIndex[4:0] ? depths_28 : _GEN_114; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_116 = 5'h1d == characterIndex[4:0] ? depths_29 : _GEN_115; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_117 = 5'h1e == characterIndex[4:0] ? depths_30 : _GEN_116; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_118 = 5'h1f == characterIndex[4:0] ? depths_31 : _GEN_117; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_120 = 5'h1 == _T_12[4:0] ? depths_1 : depths_0; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_121 = 5'h2 == _T_12[4:0] ? depths_2 : _GEN_120; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_122 = 5'h3 == _T_12[4:0] ? depths_3 : _GEN_121; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_123 = 5'h4 == _T_12[4:0] ? depths_4 : _GEN_122; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_124 = 5'h5 == _T_12[4:0] ? depths_5 : _GEN_123; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_125 = 5'h6 == _T_12[4:0] ? depths_6 : _GEN_124; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_126 = 5'h7 == _T_12[4:0] ? depths_7 : _GEN_125; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_127 = 5'h8 == _T_12[4:0] ? depths_8 : _GEN_126; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_128 = 5'h9 == _T_12[4:0] ? depths_9 : _GEN_127; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_129 = 5'ha == _T_12[4:0] ? depths_10 : _GEN_128; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_130 = 5'hb == _T_12[4:0] ? depths_11 : _GEN_129; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_131 = 5'hc == _T_12[4:0] ? depths_12 : _GEN_130; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_132 = 5'hd == _T_12[4:0] ? depths_13 : _GEN_131; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_133 = 5'he == _T_12[4:0] ? depths_14 : _GEN_132; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_134 = 5'hf == _T_12[4:0] ? depths_15 : _GEN_133; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_135 = 5'h10 == _T_12[4:0] ? depths_16 : _GEN_134; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_136 = 5'h11 == _T_12[4:0] ? depths_17 : _GEN_135; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_137 = 5'h12 == _T_12[4:0] ? depths_18 : _GEN_136; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_138 = 5'h13 == _T_12[4:0] ? depths_19 : _GEN_137; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_139 = 5'h14 == _T_12[4:0] ? depths_20 : _GEN_138; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_140 = 5'h15 == _T_12[4:0] ? depths_21 : _GEN_139; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_141 = 5'h16 == _T_12[4:0] ? depths_22 : _GEN_140; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_142 = 5'h17 == _T_12[4:0] ? depths_23 : _GEN_141; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_143 = 5'h18 == _T_12[4:0] ? depths_24 : _GEN_142; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_144 = 5'h19 == _T_12[4:0] ? depths_25 : _GEN_143; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_145 = 5'h1a == _T_12[4:0] ? depths_26 : _GEN_144; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_146 = 5'h1b == _T_12[4:0] ? depths_27 : _GEN_145; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_147 = 5'h1c == _T_12[4:0] ? depths_28 : _GEN_146; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_148 = 5'h1d == _T_12[4:0] ? depths_29 : _GEN_147; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_149 = 5'h1e == _T_12[4:0] ? depths_30 : _GEN_148; // @[codewordGenerator.scala 79:35]
  wire [3:0] _GEN_150 = 5'h1f == _T_12[4:0] ? depths_31 : _GEN_149; // @[codewordGenerator.scala 79:35]
  wire  _T_14 = _GEN_118 == _GEN_150; // @[codewordGenerator.scala 79:35]
  wire [8:0] _GEN_152 = 5'h1 == characterIndex[4:0] ? charactersIn_1 : charactersIn_0; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_153 = 5'h2 == characterIndex[4:0] ? charactersIn_2 : _GEN_152; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_154 = 5'h3 == characterIndex[4:0] ? charactersIn_3 : _GEN_153; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_155 = 5'h4 == characterIndex[4:0] ? charactersIn_4 : _GEN_154; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_156 = 5'h5 == characterIndex[4:0] ? charactersIn_5 : _GEN_155; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_157 = 5'h6 == characterIndex[4:0] ? charactersIn_6 : _GEN_156; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_158 = 5'h7 == characterIndex[4:0] ? charactersIn_7 : _GEN_157; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_159 = 5'h8 == characterIndex[4:0] ? charactersIn_8 : _GEN_158; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_160 = 5'h9 == characterIndex[4:0] ? charactersIn_9 : _GEN_159; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_161 = 5'ha == characterIndex[4:0] ? charactersIn_10 : _GEN_160; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_162 = 5'hb == characterIndex[4:0] ? charactersIn_11 : _GEN_161; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_163 = 5'hc == characterIndex[4:0] ? charactersIn_12 : _GEN_162; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_164 = 5'hd == characterIndex[4:0] ? charactersIn_13 : _GEN_163; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_165 = 5'he == characterIndex[4:0] ? charactersIn_14 : _GEN_164; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_166 = 5'hf == characterIndex[4:0] ? charactersIn_15 : _GEN_165; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_167 = 5'h10 == characterIndex[4:0] ? charactersIn_16 : _GEN_166; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_168 = 5'h11 == characterIndex[4:0] ? charactersIn_17 : _GEN_167; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_169 = 5'h12 == characterIndex[4:0] ? charactersIn_18 : _GEN_168; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_170 = 5'h13 == characterIndex[4:0] ? charactersIn_19 : _GEN_169; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_171 = 5'h14 == characterIndex[4:0] ? charactersIn_20 : _GEN_170; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_172 = 5'h15 == characterIndex[4:0] ? charactersIn_21 : _GEN_171; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_173 = 5'h16 == characterIndex[4:0] ? charactersIn_22 : _GEN_172; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_174 = 5'h17 == characterIndex[4:0] ? charactersIn_23 : _GEN_173; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_175 = 5'h18 == characterIndex[4:0] ? charactersIn_24 : _GEN_174; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_176 = 5'h19 == characterIndex[4:0] ? charactersIn_25 : _GEN_175; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_177 = 5'h1a == characterIndex[4:0] ? charactersIn_26 : _GEN_176; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_178 = 5'h1b == characterIndex[4:0] ? charactersIn_27 : _GEN_177; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_179 = 5'h1c == characterIndex[4:0] ? charactersIn_28 : _GEN_178; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_180 = 5'h1d == characterIndex[4:0] ? charactersIn_29 : _GEN_179; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_181 = 5'h1e == characterIndex[4:0] ? charactersIn_30 : _GEN_180; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_182 = 5'h1f == characterIndex[4:0] ? charactersIn_31 : _GEN_181; // @[codewordGenerator.scala 80:43]
  wire  _T_16 = _GEN_182 == 9'h100; // @[codewordGenerator.scala 80:43]
  wire [8:0] _GEN_216 = 5'h1 == _T_12[4:0] ? charactersIn_1 : charactersIn_0; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_217 = 5'h2 == _T_12[4:0] ? charactersIn_2 : _GEN_216; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_218 = 5'h3 == _T_12[4:0] ? charactersIn_3 : _GEN_217; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_219 = 5'h4 == _T_12[4:0] ? charactersIn_4 : _GEN_218; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_220 = 5'h5 == _T_12[4:0] ? charactersIn_5 : _GEN_219; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_221 = 5'h6 == _T_12[4:0] ? charactersIn_6 : _GEN_220; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_222 = 5'h7 == _T_12[4:0] ? charactersIn_7 : _GEN_221; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_223 = 5'h8 == _T_12[4:0] ? charactersIn_8 : _GEN_222; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_224 = 5'h9 == _T_12[4:0] ? charactersIn_9 : _GEN_223; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_225 = 5'ha == _T_12[4:0] ? charactersIn_10 : _GEN_224; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_226 = 5'hb == _T_12[4:0] ? charactersIn_11 : _GEN_225; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_227 = 5'hc == _T_12[4:0] ? charactersIn_12 : _GEN_226; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_228 = 5'hd == _T_12[4:0] ? charactersIn_13 : _GEN_227; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_229 = 5'he == _T_12[4:0] ? charactersIn_14 : _GEN_228; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_230 = 5'hf == _T_12[4:0] ? charactersIn_15 : _GEN_229; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_231 = 5'h10 == _T_12[4:0] ? charactersIn_16 : _GEN_230; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_232 = 5'h11 == _T_12[4:0] ? charactersIn_17 : _GEN_231; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_233 = 5'h12 == _T_12[4:0] ? charactersIn_18 : _GEN_232; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_234 = 5'h13 == _T_12[4:0] ? charactersIn_19 : _GEN_233; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_235 = 5'h14 == _T_12[4:0] ? charactersIn_20 : _GEN_234; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_236 = 5'h15 == _T_12[4:0] ? charactersIn_21 : _GEN_235; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_237 = 5'h16 == _T_12[4:0] ? charactersIn_22 : _GEN_236; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_238 = 5'h17 == _T_12[4:0] ? charactersIn_23 : _GEN_237; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_239 = 5'h18 == _T_12[4:0] ? charactersIn_24 : _GEN_238; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_240 = 5'h19 == _T_12[4:0] ? charactersIn_25 : _GEN_239; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_241 = 5'h1a == _T_12[4:0] ? charactersIn_26 : _GEN_240; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_242 = 5'h1b == _T_12[4:0] ? charactersIn_27 : _GEN_241; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_243 = 5'h1c == _T_12[4:0] ? charactersIn_28 : _GEN_242; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_244 = 5'h1d == _T_12[4:0] ? charactersIn_29 : _GEN_243; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_245 = 5'h1e == _T_12[4:0] ? charactersIn_30 : _GEN_244; // @[codewordGenerator.scala 83:40]
  wire [8:0] _GEN_246 = 5'h1f == _T_12[4:0] ? charactersIn_31 : _GEN_245; // @[codewordGenerator.scala 83:40]
  wire [8:0] _T_28 = nodes - 9'h1; // @[codewordGenerator.scala 89:36]
  wire [8:0] _GEN_9120 = {{1'd0}, characterIndex}; // @[codewordGenerator.scala 89:27]
  wire  _T_29 = _GEN_9120 >= _T_28; // @[codewordGenerator.scala 89:27]
  wire  _T_30 = state == 2'h2; // @[codewordGenerator.scala 94:21]
  wire  _T_35 = characterDepth < _GEN_118; // @[codewordGenerator.scala 99:27]
  wire [3:0] _T_39 = _GEN_118 - characterDepth; // @[codewordGenerator.scala 102:57]
  wire [30:0] _GEN_9121 = {{15'd0}, codeword}; // @[codewordGenerator.scala 102:30]
  wire [30:0] _T_40 = _GEN_9121 << _T_39; // @[codewordGenerator.scala 102:30]
  wire [15:0] _T_47 = 16'h1 << characterDepth; // @[codewordGenerator.scala 108:33]
  wire [15:0] _T_49 = _T_47 - 16'h1; // @[codewordGenerator.scala 108:52]
  wire  _T_50 = codeword != _T_49; // @[codewordGenerator.scala 108:23]
  wire [15:0] _T_52 = codeword + 16'h1; // @[codewordGenerator.scala 111:32]
  wire [15:0] _GEN_634 = _T_50 ? _T_52 : codeword; // @[codewordGenerator.scala 108:60]
  wire [4:0] _lengths_T_59 = {{1'd0}, characterDepth}; // @[codewordGenerator.scala 120:49 codewordGenerator.scala 120:49]
  wire [30:0] _GEN_1759 = _T_35 ? _T_40 : {{15'd0}, _GEN_634}; // @[codewordGenerator.scala 99:53]
  wire  _T_65 = characterIndex >= 8'hff; // @[codewordGenerator.scala 136:27]
  wire [4:0] _GEN_2296 = 8'h1 == characterIndex ? lengths_1 : lengths_0; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2297 = 8'h2 == characterIndex ? lengths_2 : _GEN_2296; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2298 = 8'h3 == characterIndex ? lengths_3 : _GEN_2297; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2299 = 8'h4 == characterIndex ? lengths_4 : _GEN_2298; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2300 = 8'h5 == characterIndex ? lengths_5 : _GEN_2299; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2301 = 8'h6 == characterIndex ? lengths_6 : _GEN_2300; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2302 = 8'h7 == characterIndex ? lengths_7 : _GEN_2301; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2303 = 8'h8 == characterIndex ? lengths_8 : _GEN_2302; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2304 = 8'h9 == characterIndex ? lengths_9 : _GEN_2303; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2305 = 8'ha == characterIndex ? lengths_10 : _GEN_2304; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2306 = 8'hb == characterIndex ? lengths_11 : _GEN_2305; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2307 = 8'hc == characterIndex ? lengths_12 : _GEN_2306; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2308 = 8'hd == characterIndex ? lengths_13 : _GEN_2307; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2309 = 8'he == characterIndex ? lengths_14 : _GEN_2308; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2310 = 8'hf == characterIndex ? lengths_15 : _GEN_2309; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2311 = 8'h10 == characterIndex ? lengths_16 : _GEN_2310; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2312 = 8'h11 == characterIndex ? lengths_17 : _GEN_2311; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2313 = 8'h12 == characterIndex ? lengths_18 : _GEN_2312; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2314 = 8'h13 == characterIndex ? lengths_19 : _GEN_2313; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2315 = 8'h14 == characterIndex ? lengths_20 : _GEN_2314; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2316 = 8'h15 == characterIndex ? lengths_21 : _GEN_2315; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2317 = 8'h16 == characterIndex ? lengths_22 : _GEN_2316; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2318 = 8'h17 == characterIndex ? lengths_23 : _GEN_2317; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2319 = 8'h18 == characterIndex ? lengths_24 : _GEN_2318; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2320 = 8'h19 == characterIndex ? lengths_25 : _GEN_2319; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2321 = 8'h1a == characterIndex ? lengths_26 : _GEN_2320; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2322 = 8'h1b == characterIndex ? lengths_27 : _GEN_2321; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2323 = 8'h1c == characterIndex ? lengths_28 : _GEN_2322; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2324 = 8'h1d == characterIndex ? lengths_29 : _GEN_2323; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2325 = 8'h1e == characterIndex ? lengths_30 : _GEN_2324; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2326 = 8'h1f == characterIndex ? lengths_31 : _GEN_2325; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2327 = 8'h20 == characterIndex ? lengths_32 : _GEN_2326; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2328 = 8'h21 == characterIndex ? lengths_33 : _GEN_2327; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2329 = 8'h22 == characterIndex ? lengths_34 : _GEN_2328; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2330 = 8'h23 == characterIndex ? lengths_35 : _GEN_2329; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2331 = 8'h24 == characterIndex ? lengths_36 : _GEN_2330; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2332 = 8'h25 == characterIndex ? lengths_37 : _GEN_2331; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2333 = 8'h26 == characterIndex ? lengths_38 : _GEN_2332; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2334 = 8'h27 == characterIndex ? lengths_39 : _GEN_2333; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2335 = 8'h28 == characterIndex ? lengths_40 : _GEN_2334; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2336 = 8'h29 == characterIndex ? lengths_41 : _GEN_2335; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2337 = 8'h2a == characterIndex ? lengths_42 : _GEN_2336; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2338 = 8'h2b == characterIndex ? lengths_43 : _GEN_2337; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2339 = 8'h2c == characterIndex ? lengths_44 : _GEN_2338; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2340 = 8'h2d == characterIndex ? lengths_45 : _GEN_2339; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2341 = 8'h2e == characterIndex ? lengths_46 : _GEN_2340; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2342 = 8'h2f == characterIndex ? lengths_47 : _GEN_2341; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2343 = 8'h30 == characterIndex ? lengths_48 : _GEN_2342; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2344 = 8'h31 == characterIndex ? lengths_49 : _GEN_2343; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2345 = 8'h32 == characterIndex ? lengths_50 : _GEN_2344; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2346 = 8'h33 == characterIndex ? lengths_51 : _GEN_2345; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2347 = 8'h34 == characterIndex ? lengths_52 : _GEN_2346; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2348 = 8'h35 == characterIndex ? lengths_53 : _GEN_2347; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2349 = 8'h36 == characterIndex ? lengths_54 : _GEN_2348; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2350 = 8'h37 == characterIndex ? lengths_55 : _GEN_2349; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2351 = 8'h38 == characterIndex ? lengths_56 : _GEN_2350; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2352 = 8'h39 == characterIndex ? lengths_57 : _GEN_2351; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2353 = 8'h3a == characterIndex ? lengths_58 : _GEN_2352; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2354 = 8'h3b == characterIndex ? lengths_59 : _GEN_2353; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2355 = 8'h3c == characterIndex ? lengths_60 : _GEN_2354; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2356 = 8'h3d == characterIndex ? lengths_61 : _GEN_2355; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2357 = 8'h3e == characterIndex ? lengths_62 : _GEN_2356; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2358 = 8'h3f == characterIndex ? lengths_63 : _GEN_2357; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2359 = 8'h40 == characterIndex ? lengths_64 : _GEN_2358; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2360 = 8'h41 == characterIndex ? lengths_65 : _GEN_2359; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2361 = 8'h42 == characterIndex ? lengths_66 : _GEN_2360; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2362 = 8'h43 == characterIndex ? lengths_67 : _GEN_2361; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2363 = 8'h44 == characterIndex ? lengths_68 : _GEN_2362; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2364 = 8'h45 == characterIndex ? lengths_69 : _GEN_2363; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2365 = 8'h46 == characterIndex ? lengths_70 : _GEN_2364; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2366 = 8'h47 == characterIndex ? lengths_71 : _GEN_2365; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2367 = 8'h48 == characterIndex ? lengths_72 : _GEN_2366; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2368 = 8'h49 == characterIndex ? lengths_73 : _GEN_2367; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2369 = 8'h4a == characterIndex ? lengths_74 : _GEN_2368; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2370 = 8'h4b == characterIndex ? lengths_75 : _GEN_2369; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2371 = 8'h4c == characterIndex ? lengths_76 : _GEN_2370; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2372 = 8'h4d == characterIndex ? lengths_77 : _GEN_2371; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2373 = 8'h4e == characterIndex ? lengths_78 : _GEN_2372; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2374 = 8'h4f == characterIndex ? lengths_79 : _GEN_2373; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2375 = 8'h50 == characterIndex ? lengths_80 : _GEN_2374; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2376 = 8'h51 == characterIndex ? lengths_81 : _GEN_2375; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2377 = 8'h52 == characterIndex ? lengths_82 : _GEN_2376; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2378 = 8'h53 == characterIndex ? lengths_83 : _GEN_2377; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2379 = 8'h54 == characterIndex ? lengths_84 : _GEN_2378; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2380 = 8'h55 == characterIndex ? lengths_85 : _GEN_2379; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2381 = 8'h56 == characterIndex ? lengths_86 : _GEN_2380; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2382 = 8'h57 == characterIndex ? lengths_87 : _GEN_2381; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2383 = 8'h58 == characterIndex ? lengths_88 : _GEN_2382; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2384 = 8'h59 == characterIndex ? lengths_89 : _GEN_2383; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2385 = 8'h5a == characterIndex ? lengths_90 : _GEN_2384; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2386 = 8'h5b == characterIndex ? lengths_91 : _GEN_2385; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2387 = 8'h5c == characterIndex ? lengths_92 : _GEN_2386; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2388 = 8'h5d == characterIndex ? lengths_93 : _GEN_2387; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2389 = 8'h5e == characterIndex ? lengths_94 : _GEN_2388; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2390 = 8'h5f == characterIndex ? lengths_95 : _GEN_2389; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2391 = 8'h60 == characterIndex ? lengths_96 : _GEN_2390; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2392 = 8'h61 == characterIndex ? lengths_97 : _GEN_2391; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2393 = 8'h62 == characterIndex ? lengths_98 : _GEN_2392; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2394 = 8'h63 == characterIndex ? lengths_99 : _GEN_2393; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2395 = 8'h64 == characterIndex ? lengths_100 : _GEN_2394; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2396 = 8'h65 == characterIndex ? lengths_101 : _GEN_2395; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2397 = 8'h66 == characterIndex ? lengths_102 : _GEN_2396; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2398 = 8'h67 == characterIndex ? lengths_103 : _GEN_2397; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2399 = 8'h68 == characterIndex ? lengths_104 : _GEN_2398; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2400 = 8'h69 == characterIndex ? lengths_105 : _GEN_2399; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2401 = 8'h6a == characterIndex ? lengths_106 : _GEN_2400; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2402 = 8'h6b == characterIndex ? lengths_107 : _GEN_2401; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2403 = 8'h6c == characterIndex ? lengths_108 : _GEN_2402; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2404 = 8'h6d == characterIndex ? lengths_109 : _GEN_2403; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2405 = 8'h6e == characterIndex ? lengths_110 : _GEN_2404; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2406 = 8'h6f == characterIndex ? lengths_111 : _GEN_2405; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2407 = 8'h70 == characterIndex ? lengths_112 : _GEN_2406; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2408 = 8'h71 == characterIndex ? lengths_113 : _GEN_2407; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2409 = 8'h72 == characterIndex ? lengths_114 : _GEN_2408; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2410 = 8'h73 == characterIndex ? lengths_115 : _GEN_2409; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2411 = 8'h74 == characterIndex ? lengths_116 : _GEN_2410; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2412 = 8'h75 == characterIndex ? lengths_117 : _GEN_2411; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2413 = 8'h76 == characterIndex ? lengths_118 : _GEN_2412; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2414 = 8'h77 == characterIndex ? lengths_119 : _GEN_2413; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2415 = 8'h78 == characterIndex ? lengths_120 : _GEN_2414; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2416 = 8'h79 == characterIndex ? lengths_121 : _GEN_2415; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2417 = 8'h7a == characterIndex ? lengths_122 : _GEN_2416; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2418 = 8'h7b == characterIndex ? lengths_123 : _GEN_2417; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2419 = 8'h7c == characterIndex ? lengths_124 : _GEN_2418; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2420 = 8'h7d == characterIndex ? lengths_125 : _GEN_2419; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2421 = 8'h7e == characterIndex ? lengths_126 : _GEN_2420; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2422 = 8'h7f == characterIndex ? lengths_127 : _GEN_2421; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2423 = 8'h80 == characterIndex ? lengths_128 : _GEN_2422; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2424 = 8'h81 == characterIndex ? lengths_129 : _GEN_2423; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2425 = 8'h82 == characterIndex ? lengths_130 : _GEN_2424; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2426 = 8'h83 == characterIndex ? lengths_131 : _GEN_2425; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2427 = 8'h84 == characterIndex ? lengths_132 : _GEN_2426; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2428 = 8'h85 == characterIndex ? lengths_133 : _GEN_2427; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2429 = 8'h86 == characterIndex ? lengths_134 : _GEN_2428; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2430 = 8'h87 == characterIndex ? lengths_135 : _GEN_2429; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2431 = 8'h88 == characterIndex ? lengths_136 : _GEN_2430; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2432 = 8'h89 == characterIndex ? lengths_137 : _GEN_2431; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2433 = 8'h8a == characterIndex ? lengths_138 : _GEN_2432; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2434 = 8'h8b == characterIndex ? lengths_139 : _GEN_2433; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2435 = 8'h8c == characterIndex ? lengths_140 : _GEN_2434; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2436 = 8'h8d == characterIndex ? lengths_141 : _GEN_2435; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2437 = 8'h8e == characterIndex ? lengths_142 : _GEN_2436; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2438 = 8'h8f == characterIndex ? lengths_143 : _GEN_2437; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2439 = 8'h90 == characterIndex ? lengths_144 : _GEN_2438; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2440 = 8'h91 == characterIndex ? lengths_145 : _GEN_2439; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2441 = 8'h92 == characterIndex ? lengths_146 : _GEN_2440; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2442 = 8'h93 == characterIndex ? lengths_147 : _GEN_2441; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2443 = 8'h94 == characterIndex ? lengths_148 : _GEN_2442; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2444 = 8'h95 == characterIndex ? lengths_149 : _GEN_2443; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2445 = 8'h96 == characterIndex ? lengths_150 : _GEN_2444; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2446 = 8'h97 == characterIndex ? lengths_151 : _GEN_2445; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2447 = 8'h98 == characterIndex ? lengths_152 : _GEN_2446; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2448 = 8'h99 == characterIndex ? lengths_153 : _GEN_2447; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2449 = 8'h9a == characterIndex ? lengths_154 : _GEN_2448; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2450 = 8'h9b == characterIndex ? lengths_155 : _GEN_2449; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2451 = 8'h9c == characterIndex ? lengths_156 : _GEN_2450; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2452 = 8'h9d == characterIndex ? lengths_157 : _GEN_2451; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2453 = 8'h9e == characterIndex ? lengths_158 : _GEN_2452; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2454 = 8'h9f == characterIndex ? lengths_159 : _GEN_2453; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2455 = 8'ha0 == characterIndex ? lengths_160 : _GEN_2454; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2456 = 8'ha1 == characterIndex ? lengths_161 : _GEN_2455; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2457 = 8'ha2 == characterIndex ? lengths_162 : _GEN_2456; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2458 = 8'ha3 == characterIndex ? lengths_163 : _GEN_2457; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2459 = 8'ha4 == characterIndex ? lengths_164 : _GEN_2458; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2460 = 8'ha5 == characterIndex ? lengths_165 : _GEN_2459; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2461 = 8'ha6 == characterIndex ? lengths_166 : _GEN_2460; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2462 = 8'ha7 == characterIndex ? lengths_167 : _GEN_2461; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2463 = 8'ha8 == characterIndex ? lengths_168 : _GEN_2462; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2464 = 8'ha9 == characterIndex ? lengths_169 : _GEN_2463; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2465 = 8'haa == characterIndex ? lengths_170 : _GEN_2464; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2466 = 8'hab == characterIndex ? lengths_171 : _GEN_2465; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2467 = 8'hac == characterIndex ? lengths_172 : _GEN_2466; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2468 = 8'had == characterIndex ? lengths_173 : _GEN_2467; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2469 = 8'hae == characterIndex ? lengths_174 : _GEN_2468; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2470 = 8'haf == characterIndex ? lengths_175 : _GEN_2469; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2471 = 8'hb0 == characterIndex ? lengths_176 : _GEN_2470; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2472 = 8'hb1 == characterIndex ? lengths_177 : _GEN_2471; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2473 = 8'hb2 == characterIndex ? lengths_178 : _GEN_2472; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2474 = 8'hb3 == characterIndex ? lengths_179 : _GEN_2473; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2475 = 8'hb4 == characterIndex ? lengths_180 : _GEN_2474; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2476 = 8'hb5 == characterIndex ? lengths_181 : _GEN_2475; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2477 = 8'hb6 == characterIndex ? lengths_182 : _GEN_2476; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2478 = 8'hb7 == characterIndex ? lengths_183 : _GEN_2477; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2479 = 8'hb8 == characterIndex ? lengths_184 : _GEN_2478; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2480 = 8'hb9 == characterIndex ? lengths_185 : _GEN_2479; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2481 = 8'hba == characterIndex ? lengths_186 : _GEN_2480; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2482 = 8'hbb == characterIndex ? lengths_187 : _GEN_2481; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2483 = 8'hbc == characterIndex ? lengths_188 : _GEN_2482; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2484 = 8'hbd == characterIndex ? lengths_189 : _GEN_2483; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2485 = 8'hbe == characterIndex ? lengths_190 : _GEN_2484; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2486 = 8'hbf == characterIndex ? lengths_191 : _GEN_2485; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2487 = 8'hc0 == characterIndex ? lengths_192 : _GEN_2486; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2488 = 8'hc1 == characterIndex ? lengths_193 : _GEN_2487; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2489 = 8'hc2 == characterIndex ? lengths_194 : _GEN_2488; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2490 = 8'hc3 == characterIndex ? lengths_195 : _GEN_2489; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2491 = 8'hc4 == characterIndex ? lengths_196 : _GEN_2490; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2492 = 8'hc5 == characterIndex ? lengths_197 : _GEN_2491; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2493 = 8'hc6 == characterIndex ? lengths_198 : _GEN_2492; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2494 = 8'hc7 == characterIndex ? lengths_199 : _GEN_2493; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2495 = 8'hc8 == characterIndex ? lengths_200 : _GEN_2494; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2496 = 8'hc9 == characterIndex ? lengths_201 : _GEN_2495; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2497 = 8'hca == characterIndex ? lengths_202 : _GEN_2496; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2498 = 8'hcb == characterIndex ? lengths_203 : _GEN_2497; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2499 = 8'hcc == characterIndex ? lengths_204 : _GEN_2498; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2500 = 8'hcd == characterIndex ? lengths_205 : _GEN_2499; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2501 = 8'hce == characterIndex ? lengths_206 : _GEN_2500; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2502 = 8'hcf == characterIndex ? lengths_207 : _GEN_2501; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2503 = 8'hd0 == characterIndex ? lengths_208 : _GEN_2502; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2504 = 8'hd1 == characterIndex ? lengths_209 : _GEN_2503; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2505 = 8'hd2 == characterIndex ? lengths_210 : _GEN_2504; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2506 = 8'hd3 == characterIndex ? lengths_211 : _GEN_2505; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2507 = 8'hd4 == characterIndex ? lengths_212 : _GEN_2506; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2508 = 8'hd5 == characterIndex ? lengths_213 : _GEN_2507; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2509 = 8'hd6 == characterIndex ? lengths_214 : _GEN_2508; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2510 = 8'hd7 == characterIndex ? lengths_215 : _GEN_2509; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2511 = 8'hd8 == characterIndex ? lengths_216 : _GEN_2510; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2512 = 8'hd9 == characterIndex ? lengths_217 : _GEN_2511; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2513 = 8'hda == characterIndex ? lengths_218 : _GEN_2512; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2514 = 8'hdb == characterIndex ? lengths_219 : _GEN_2513; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2515 = 8'hdc == characterIndex ? lengths_220 : _GEN_2514; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2516 = 8'hdd == characterIndex ? lengths_221 : _GEN_2515; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2517 = 8'hde == characterIndex ? lengths_222 : _GEN_2516; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2518 = 8'hdf == characterIndex ? lengths_223 : _GEN_2517; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2519 = 8'he0 == characterIndex ? lengths_224 : _GEN_2518; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2520 = 8'he1 == characterIndex ? lengths_225 : _GEN_2519; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2521 = 8'he2 == characterIndex ? lengths_226 : _GEN_2520; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2522 = 8'he3 == characterIndex ? lengths_227 : _GEN_2521; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2523 = 8'he4 == characterIndex ? lengths_228 : _GEN_2522; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2524 = 8'he5 == characterIndex ? lengths_229 : _GEN_2523; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2525 = 8'he6 == characterIndex ? lengths_230 : _GEN_2524; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2526 = 8'he7 == characterIndex ? lengths_231 : _GEN_2525; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2527 = 8'he8 == characterIndex ? lengths_232 : _GEN_2526; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2528 = 8'he9 == characterIndex ? lengths_233 : _GEN_2527; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2529 = 8'hea == characterIndex ? lengths_234 : _GEN_2528; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2530 = 8'heb == characterIndex ? lengths_235 : _GEN_2529; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2531 = 8'hec == characterIndex ? lengths_236 : _GEN_2530; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2532 = 8'hed == characterIndex ? lengths_237 : _GEN_2531; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2533 = 8'hee == characterIndex ? lengths_238 : _GEN_2532; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2534 = 8'hef == characterIndex ? lengths_239 : _GEN_2533; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2535 = 8'hf0 == characterIndex ? lengths_240 : _GEN_2534; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2536 = 8'hf1 == characterIndex ? lengths_241 : _GEN_2535; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2537 = 8'hf2 == characterIndex ? lengths_242 : _GEN_2536; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2538 = 8'hf3 == characterIndex ? lengths_243 : _GEN_2537; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2539 = 8'hf4 == characterIndex ? lengths_244 : _GEN_2538; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2540 = 8'hf5 == characterIndex ? lengths_245 : _GEN_2539; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2541 = 8'hf6 == characterIndex ? lengths_246 : _GEN_2540; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2542 = 8'hf7 == characterIndex ? lengths_247 : _GEN_2541; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2543 = 8'hf8 == characterIndex ? lengths_248 : _GEN_2542; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2544 = 8'hf9 == characterIndex ? lengths_249 : _GEN_2543; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2545 = 8'hfa == characterIndex ? lengths_250 : _GEN_2544; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2546 = 8'hfb == characterIndex ? lengths_251 : _GEN_2545; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2547 = 8'hfc == characterIndex ? lengths_252 : _GEN_2546; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2548 = 8'hfd == characterIndex ? lengths_253 : _GEN_2547; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2549 = 8'hfe == characterIndex ? lengths_254 : _GEN_2548; // @[codewordGenerator.scala 139:36]
  wire [4:0] _GEN_2550 = 8'hff == characterIndex ? lengths_255 : _GEN_2549; // @[codewordGenerator.scala 139:36]
  wire  _T_66 = _GEN_2550 == 5'h0; // @[codewordGenerator.scala 139:36]
  wire [23:0] _T_67 = {escapeCodeword,characterIndex}; // @[Cat.scala 29:58]
  wire [4:0] _GEN_9123 = {{1'd0}, escapeCharacterLength}; // @[codewordGenerator.scala 142:61]
  wire [4:0] _T_69 = _GEN_9123 + 5'h8; // @[codewordGenerator.scala 142:61]
  wire [15:0] _GEN_3576 = 8'h1 == characterIndex ? codewords_1 : codewords_0; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3577 = 8'h2 == characterIndex ? codewords_2 : _GEN_3576; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3578 = 8'h3 == characterIndex ? codewords_3 : _GEN_3577; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3579 = 8'h4 == characterIndex ? codewords_4 : _GEN_3578; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3580 = 8'h5 == characterIndex ? codewords_5 : _GEN_3579; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3581 = 8'h6 == characterIndex ? codewords_6 : _GEN_3580; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3582 = 8'h7 == characterIndex ? codewords_7 : _GEN_3581; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3583 = 8'h8 == characterIndex ? codewords_8 : _GEN_3582; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3584 = 8'h9 == characterIndex ? codewords_9 : _GEN_3583; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3585 = 8'ha == characterIndex ? codewords_10 : _GEN_3584; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3586 = 8'hb == characterIndex ? codewords_11 : _GEN_3585; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3587 = 8'hc == characterIndex ? codewords_12 : _GEN_3586; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3588 = 8'hd == characterIndex ? codewords_13 : _GEN_3587; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3589 = 8'he == characterIndex ? codewords_14 : _GEN_3588; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3590 = 8'hf == characterIndex ? codewords_15 : _GEN_3589; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3591 = 8'h10 == characterIndex ? codewords_16 : _GEN_3590; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3592 = 8'h11 == characterIndex ? codewords_17 : _GEN_3591; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3593 = 8'h12 == characterIndex ? codewords_18 : _GEN_3592; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3594 = 8'h13 == characterIndex ? codewords_19 : _GEN_3593; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3595 = 8'h14 == characterIndex ? codewords_20 : _GEN_3594; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3596 = 8'h15 == characterIndex ? codewords_21 : _GEN_3595; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3597 = 8'h16 == characterIndex ? codewords_22 : _GEN_3596; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3598 = 8'h17 == characterIndex ? codewords_23 : _GEN_3597; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3599 = 8'h18 == characterIndex ? codewords_24 : _GEN_3598; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3600 = 8'h19 == characterIndex ? codewords_25 : _GEN_3599; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3601 = 8'h1a == characterIndex ? codewords_26 : _GEN_3600; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3602 = 8'h1b == characterIndex ? codewords_27 : _GEN_3601; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3603 = 8'h1c == characterIndex ? codewords_28 : _GEN_3602; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3604 = 8'h1d == characterIndex ? codewords_29 : _GEN_3603; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3605 = 8'h1e == characterIndex ? codewords_30 : _GEN_3604; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3606 = 8'h1f == characterIndex ? codewords_31 : _GEN_3605; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3607 = 8'h20 == characterIndex ? codewords_32 : _GEN_3606; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3608 = 8'h21 == characterIndex ? codewords_33 : _GEN_3607; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3609 = 8'h22 == characterIndex ? codewords_34 : _GEN_3608; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3610 = 8'h23 == characterIndex ? codewords_35 : _GEN_3609; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3611 = 8'h24 == characterIndex ? codewords_36 : _GEN_3610; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3612 = 8'h25 == characterIndex ? codewords_37 : _GEN_3611; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3613 = 8'h26 == characterIndex ? codewords_38 : _GEN_3612; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3614 = 8'h27 == characterIndex ? codewords_39 : _GEN_3613; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3615 = 8'h28 == characterIndex ? codewords_40 : _GEN_3614; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3616 = 8'h29 == characterIndex ? codewords_41 : _GEN_3615; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3617 = 8'h2a == characterIndex ? codewords_42 : _GEN_3616; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3618 = 8'h2b == characterIndex ? codewords_43 : _GEN_3617; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3619 = 8'h2c == characterIndex ? codewords_44 : _GEN_3618; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3620 = 8'h2d == characterIndex ? codewords_45 : _GEN_3619; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3621 = 8'h2e == characterIndex ? codewords_46 : _GEN_3620; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3622 = 8'h2f == characterIndex ? codewords_47 : _GEN_3621; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3623 = 8'h30 == characterIndex ? codewords_48 : _GEN_3622; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3624 = 8'h31 == characterIndex ? codewords_49 : _GEN_3623; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3625 = 8'h32 == characterIndex ? codewords_50 : _GEN_3624; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3626 = 8'h33 == characterIndex ? codewords_51 : _GEN_3625; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3627 = 8'h34 == characterIndex ? codewords_52 : _GEN_3626; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3628 = 8'h35 == characterIndex ? codewords_53 : _GEN_3627; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3629 = 8'h36 == characterIndex ? codewords_54 : _GEN_3628; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3630 = 8'h37 == characterIndex ? codewords_55 : _GEN_3629; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3631 = 8'h38 == characterIndex ? codewords_56 : _GEN_3630; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3632 = 8'h39 == characterIndex ? codewords_57 : _GEN_3631; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3633 = 8'h3a == characterIndex ? codewords_58 : _GEN_3632; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3634 = 8'h3b == characterIndex ? codewords_59 : _GEN_3633; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3635 = 8'h3c == characterIndex ? codewords_60 : _GEN_3634; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3636 = 8'h3d == characterIndex ? codewords_61 : _GEN_3635; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3637 = 8'h3e == characterIndex ? codewords_62 : _GEN_3636; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3638 = 8'h3f == characterIndex ? codewords_63 : _GEN_3637; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3639 = 8'h40 == characterIndex ? codewords_64 : _GEN_3638; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3640 = 8'h41 == characterIndex ? codewords_65 : _GEN_3639; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3641 = 8'h42 == characterIndex ? codewords_66 : _GEN_3640; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3642 = 8'h43 == characterIndex ? codewords_67 : _GEN_3641; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3643 = 8'h44 == characterIndex ? codewords_68 : _GEN_3642; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3644 = 8'h45 == characterIndex ? codewords_69 : _GEN_3643; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3645 = 8'h46 == characterIndex ? codewords_70 : _GEN_3644; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3646 = 8'h47 == characterIndex ? codewords_71 : _GEN_3645; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3647 = 8'h48 == characterIndex ? codewords_72 : _GEN_3646; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3648 = 8'h49 == characterIndex ? codewords_73 : _GEN_3647; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3649 = 8'h4a == characterIndex ? codewords_74 : _GEN_3648; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3650 = 8'h4b == characterIndex ? codewords_75 : _GEN_3649; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3651 = 8'h4c == characterIndex ? codewords_76 : _GEN_3650; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3652 = 8'h4d == characterIndex ? codewords_77 : _GEN_3651; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3653 = 8'h4e == characterIndex ? codewords_78 : _GEN_3652; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3654 = 8'h4f == characterIndex ? codewords_79 : _GEN_3653; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3655 = 8'h50 == characterIndex ? codewords_80 : _GEN_3654; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3656 = 8'h51 == characterIndex ? codewords_81 : _GEN_3655; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3657 = 8'h52 == characterIndex ? codewords_82 : _GEN_3656; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3658 = 8'h53 == characterIndex ? codewords_83 : _GEN_3657; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3659 = 8'h54 == characterIndex ? codewords_84 : _GEN_3658; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3660 = 8'h55 == characterIndex ? codewords_85 : _GEN_3659; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3661 = 8'h56 == characterIndex ? codewords_86 : _GEN_3660; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3662 = 8'h57 == characterIndex ? codewords_87 : _GEN_3661; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3663 = 8'h58 == characterIndex ? codewords_88 : _GEN_3662; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3664 = 8'h59 == characterIndex ? codewords_89 : _GEN_3663; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3665 = 8'h5a == characterIndex ? codewords_90 : _GEN_3664; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3666 = 8'h5b == characterIndex ? codewords_91 : _GEN_3665; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3667 = 8'h5c == characterIndex ? codewords_92 : _GEN_3666; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3668 = 8'h5d == characterIndex ? codewords_93 : _GEN_3667; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3669 = 8'h5e == characterIndex ? codewords_94 : _GEN_3668; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3670 = 8'h5f == characterIndex ? codewords_95 : _GEN_3669; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3671 = 8'h60 == characterIndex ? codewords_96 : _GEN_3670; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3672 = 8'h61 == characterIndex ? codewords_97 : _GEN_3671; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3673 = 8'h62 == characterIndex ? codewords_98 : _GEN_3672; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3674 = 8'h63 == characterIndex ? codewords_99 : _GEN_3673; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3675 = 8'h64 == characterIndex ? codewords_100 : _GEN_3674; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3676 = 8'h65 == characterIndex ? codewords_101 : _GEN_3675; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3677 = 8'h66 == characterIndex ? codewords_102 : _GEN_3676; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3678 = 8'h67 == characterIndex ? codewords_103 : _GEN_3677; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3679 = 8'h68 == characterIndex ? codewords_104 : _GEN_3678; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3680 = 8'h69 == characterIndex ? codewords_105 : _GEN_3679; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3681 = 8'h6a == characterIndex ? codewords_106 : _GEN_3680; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3682 = 8'h6b == characterIndex ? codewords_107 : _GEN_3681; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3683 = 8'h6c == characterIndex ? codewords_108 : _GEN_3682; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3684 = 8'h6d == characterIndex ? codewords_109 : _GEN_3683; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3685 = 8'h6e == characterIndex ? codewords_110 : _GEN_3684; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3686 = 8'h6f == characterIndex ? codewords_111 : _GEN_3685; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3687 = 8'h70 == characterIndex ? codewords_112 : _GEN_3686; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3688 = 8'h71 == characterIndex ? codewords_113 : _GEN_3687; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3689 = 8'h72 == characterIndex ? codewords_114 : _GEN_3688; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3690 = 8'h73 == characterIndex ? codewords_115 : _GEN_3689; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3691 = 8'h74 == characterIndex ? codewords_116 : _GEN_3690; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3692 = 8'h75 == characterIndex ? codewords_117 : _GEN_3691; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3693 = 8'h76 == characterIndex ? codewords_118 : _GEN_3692; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3694 = 8'h77 == characterIndex ? codewords_119 : _GEN_3693; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3695 = 8'h78 == characterIndex ? codewords_120 : _GEN_3694; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3696 = 8'h79 == characterIndex ? codewords_121 : _GEN_3695; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3697 = 8'h7a == characterIndex ? codewords_122 : _GEN_3696; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3698 = 8'h7b == characterIndex ? codewords_123 : _GEN_3697; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3699 = 8'h7c == characterIndex ? codewords_124 : _GEN_3698; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3700 = 8'h7d == characterIndex ? codewords_125 : _GEN_3699; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3701 = 8'h7e == characterIndex ? codewords_126 : _GEN_3700; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3702 = 8'h7f == characterIndex ? codewords_127 : _GEN_3701; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3703 = 8'h80 == characterIndex ? codewords_128 : _GEN_3702; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3704 = 8'h81 == characterIndex ? codewords_129 : _GEN_3703; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3705 = 8'h82 == characterIndex ? codewords_130 : _GEN_3704; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3706 = 8'h83 == characterIndex ? codewords_131 : _GEN_3705; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3707 = 8'h84 == characterIndex ? codewords_132 : _GEN_3706; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3708 = 8'h85 == characterIndex ? codewords_133 : _GEN_3707; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3709 = 8'h86 == characterIndex ? codewords_134 : _GEN_3708; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3710 = 8'h87 == characterIndex ? codewords_135 : _GEN_3709; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3711 = 8'h88 == characterIndex ? codewords_136 : _GEN_3710; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3712 = 8'h89 == characterIndex ? codewords_137 : _GEN_3711; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3713 = 8'h8a == characterIndex ? codewords_138 : _GEN_3712; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3714 = 8'h8b == characterIndex ? codewords_139 : _GEN_3713; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3715 = 8'h8c == characterIndex ? codewords_140 : _GEN_3714; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3716 = 8'h8d == characterIndex ? codewords_141 : _GEN_3715; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3717 = 8'h8e == characterIndex ? codewords_142 : _GEN_3716; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3718 = 8'h8f == characterIndex ? codewords_143 : _GEN_3717; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3719 = 8'h90 == characterIndex ? codewords_144 : _GEN_3718; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3720 = 8'h91 == characterIndex ? codewords_145 : _GEN_3719; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3721 = 8'h92 == characterIndex ? codewords_146 : _GEN_3720; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3722 = 8'h93 == characterIndex ? codewords_147 : _GEN_3721; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3723 = 8'h94 == characterIndex ? codewords_148 : _GEN_3722; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3724 = 8'h95 == characterIndex ? codewords_149 : _GEN_3723; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3725 = 8'h96 == characterIndex ? codewords_150 : _GEN_3724; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3726 = 8'h97 == characterIndex ? codewords_151 : _GEN_3725; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3727 = 8'h98 == characterIndex ? codewords_152 : _GEN_3726; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3728 = 8'h99 == characterIndex ? codewords_153 : _GEN_3727; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3729 = 8'h9a == characterIndex ? codewords_154 : _GEN_3728; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3730 = 8'h9b == characterIndex ? codewords_155 : _GEN_3729; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3731 = 8'h9c == characterIndex ? codewords_156 : _GEN_3730; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3732 = 8'h9d == characterIndex ? codewords_157 : _GEN_3731; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3733 = 8'h9e == characterIndex ? codewords_158 : _GEN_3732; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3734 = 8'h9f == characterIndex ? codewords_159 : _GEN_3733; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3735 = 8'ha0 == characterIndex ? codewords_160 : _GEN_3734; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3736 = 8'ha1 == characterIndex ? codewords_161 : _GEN_3735; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3737 = 8'ha2 == characterIndex ? codewords_162 : _GEN_3736; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3738 = 8'ha3 == characterIndex ? codewords_163 : _GEN_3737; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3739 = 8'ha4 == characterIndex ? codewords_164 : _GEN_3738; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3740 = 8'ha5 == characterIndex ? codewords_165 : _GEN_3739; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3741 = 8'ha6 == characterIndex ? codewords_166 : _GEN_3740; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3742 = 8'ha7 == characterIndex ? codewords_167 : _GEN_3741; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3743 = 8'ha8 == characterIndex ? codewords_168 : _GEN_3742; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3744 = 8'ha9 == characterIndex ? codewords_169 : _GEN_3743; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3745 = 8'haa == characterIndex ? codewords_170 : _GEN_3744; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3746 = 8'hab == characterIndex ? codewords_171 : _GEN_3745; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3747 = 8'hac == characterIndex ? codewords_172 : _GEN_3746; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3748 = 8'had == characterIndex ? codewords_173 : _GEN_3747; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3749 = 8'hae == characterIndex ? codewords_174 : _GEN_3748; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3750 = 8'haf == characterIndex ? codewords_175 : _GEN_3749; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3751 = 8'hb0 == characterIndex ? codewords_176 : _GEN_3750; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3752 = 8'hb1 == characterIndex ? codewords_177 : _GEN_3751; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3753 = 8'hb2 == characterIndex ? codewords_178 : _GEN_3752; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3754 = 8'hb3 == characterIndex ? codewords_179 : _GEN_3753; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3755 = 8'hb4 == characterIndex ? codewords_180 : _GEN_3754; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3756 = 8'hb5 == characterIndex ? codewords_181 : _GEN_3755; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3757 = 8'hb6 == characterIndex ? codewords_182 : _GEN_3756; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3758 = 8'hb7 == characterIndex ? codewords_183 : _GEN_3757; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3759 = 8'hb8 == characterIndex ? codewords_184 : _GEN_3758; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3760 = 8'hb9 == characterIndex ? codewords_185 : _GEN_3759; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3761 = 8'hba == characterIndex ? codewords_186 : _GEN_3760; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3762 = 8'hbb == characterIndex ? codewords_187 : _GEN_3761; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3763 = 8'hbc == characterIndex ? codewords_188 : _GEN_3762; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3764 = 8'hbd == characterIndex ? codewords_189 : _GEN_3763; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3765 = 8'hbe == characterIndex ? codewords_190 : _GEN_3764; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3766 = 8'hbf == characterIndex ? codewords_191 : _GEN_3765; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3767 = 8'hc0 == characterIndex ? codewords_192 : _GEN_3766; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3768 = 8'hc1 == characterIndex ? codewords_193 : _GEN_3767; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3769 = 8'hc2 == characterIndex ? codewords_194 : _GEN_3768; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3770 = 8'hc3 == characterIndex ? codewords_195 : _GEN_3769; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3771 = 8'hc4 == characterIndex ? codewords_196 : _GEN_3770; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3772 = 8'hc5 == characterIndex ? codewords_197 : _GEN_3771; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3773 = 8'hc6 == characterIndex ? codewords_198 : _GEN_3772; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3774 = 8'hc7 == characterIndex ? codewords_199 : _GEN_3773; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3775 = 8'hc8 == characterIndex ? codewords_200 : _GEN_3774; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3776 = 8'hc9 == characterIndex ? codewords_201 : _GEN_3775; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3777 = 8'hca == characterIndex ? codewords_202 : _GEN_3776; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3778 = 8'hcb == characterIndex ? codewords_203 : _GEN_3777; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3779 = 8'hcc == characterIndex ? codewords_204 : _GEN_3778; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3780 = 8'hcd == characterIndex ? codewords_205 : _GEN_3779; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3781 = 8'hce == characterIndex ? codewords_206 : _GEN_3780; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3782 = 8'hcf == characterIndex ? codewords_207 : _GEN_3781; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3783 = 8'hd0 == characterIndex ? codewords_208 : _GEN_3782; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3784 = 8'hd1 == characterIndex ? codewords_209 : _GEN_3783; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3785 = 8'hd2 == characterIndex ? codewords_210 : _GEN_3784; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3786 = 8'hd3 == characterIndex ? codewords_211 : _GEN_3785; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3787 = 8'hd4 == characterIndex ? codewords_212 : _GEN_3786; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3788 = 8'hd5 == characterIndex ? codewords_213 : _GEN_3787; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3789 = 8'hd6 == characterIndex ? codewords_214 : _GEN_3788; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3790 = 8'hd7 == characterIndex ? codewords_215 : _GEN_3789; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3791 = 8'hd8 == characterIndex ? codewords_216 : _GEN_3790; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3792 = 8'hd9 == characterIndex ? codewords_217 : _GEN_3791; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3793 = 8'hda == characterIndex ? codewords_218 : _GEN_3792; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3794 = 8'hdb == characterIndex ? codewords_219 : _GEN_3793; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3795 = 8'hdc == characterIndex ? codewords_220 : _GEN_3794; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3796 = 8'hdd == characterIndex ? codewords_221 : _GEN_3795; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3797 = 8'hde == characterIndex ? codewords_222 : _GEN_3796; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3798 = 8'hdf == characterIndex ? codewords_223 : _GEN_3797; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3799 = 8'he0 == characterIndex ? codewords_224 : _GEN_3798; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3800 = 8'he1 == characterIndex ? codewords_225 : _GEN_3799; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3801 = 8'he2 == characterIndex ? codewords_226 : _GEN_3800; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3802 = 8'he3 == characterIndex ? codewords_227 : _GEN_3801; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3803 = 8'he4 == characterIndex ? codewords_228 : _GEN_3802; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3804 = 8'he5 == characterIndex ? codewords_229 : _GEN_3803; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3805 = 8'he6 == characterIndex ? codewords_230 : _GEN_3804; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3806 = 8'he7 == characterIndex ? codewords_231 : _GEN_3805; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3807 = 8'he8 == characterIndex ? codewords_232 : _GEN_3806; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3808 = 8'he9 == characterIndex ? codewords_233 : _GEN_3807; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3809 = 8'hea == characterIndex ? codewords_234 : _GEN_3808; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3810 = 8'heb == characterIndex ? codewords_235 : _GEN_3809; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3811 = 8'hec == characterIndex ? codewords_236 : _GEN_3810; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3812 = 8'hed == characterIndex ? codewords_237 : _GEN_3811; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3813 = 8'hee == characterIndex ? codewords_238 : _GEN_3812; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3814 = 8'hef == characterIndex ? codewords_239 : _GEN_3813; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3815 = 8'hf0 == characterIndex ? codewords_240 : _GEN_3814; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3816 = 8'hf1 == characterIndex ? codewords_241 : _GEN_3815; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3817 = 8'hf2 == characterIndex ? codewords_242 : _GEN_3816; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3818 = 8'hf3 == characterIndex ? codewords_243 : _GEN_3817; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3819 = 8'hf4 == characterIndex ? codewords_244 : _GEN_3818; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3820 = 8'hf5 == characterIndex ? codewords_245 : _GEN_3819; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3821 = 8'hf6 == characterIndex ? codewords_246 : _GEN_3820; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3822 = 8'hf7 == characterIndex ? codewords_247 : _GEN_3821; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3823 = 8'hf8 == characterIndex ? codewords_248 : _GEN_3822; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3824 = 8'hf9 == characterIndex ? codewords_249 : _GEN_3823; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3825 = 8'hfa == characterIndex ? codewords_250 : _GEN_3824; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3826 = 8'hfb == characterIndex ? codewords_251 : _GEN_3825; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3827 = 8'hfc == characterIndex ? codewords_252 : _GEN_3826; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3828 = 8'hfd == characterIndex ? codewords_253 : _GEN_3827; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3829 = 8'hfe == characterIndex ? codewords_254 : _GEN_3828; // @[codewordGenerator.scala 145:38]
  wire [15:0] _GEN_3830 = 8'hff == characterIndex ? codewords_255 : _GEN_3829; // @[codewordGenerator.scala 145:38]
  wire [23:0] _codewordsOut_characterIndex_0 = {{8'd0}, _GEN_3830}; // @[codewordGenerator.scala 145:38 codewordGenerator.scala 145:38]
  wire [30:0] _GEN_5113 = _T_30 ? _GEN_1759 : {{15'd0}, codeword}; // @[codewordGenerator.scala 94:47]
  wire [30:0] _GEN_6451 = _T_9 ? {{15'd0}, codeword} : _GEN_5113; // @[codewordGenerator.scala 76:43]
  wire [7:0] _GEN_7784 = _T_6 ? _GEN_33 : {{4'd0}, depths_0}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7785 = _T_6 ? _GEN_34 : {{4'd0}, depths_1}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7786 = _T_6 ? _GEN_35 : {{4'd0}, depths_2}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7787 = _T_6 ? _GEN_36 : {{4'd0}, depths_3}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7788 = _T_6 ? _GEN_37 : {{4'd0}, depths_4}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7789 = _T_6 ? _GEN_38 : {{4'd0}, depths_5}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7790 = _T_6 ? _GEN_39 : {{4'd0}, depths_6}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7791 = _T_6 ? _GEN_40 : {{4'd0}, depths_7}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7792 = _T_6 ? _GEN_41 : {{4'd0}, depths_8}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7793 = _T_6 ? _GEN_42 : {{4'd0}, depths_9}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7794 = _T_6 ? _GEN_43 : {{4'd0}, depths_10}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7795 = _T_6 ? _GEN_44 : {{4'd0}, depths_11}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7796 = _T_6 ? _GEN_45 : {{4'd0}, depths_12}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7797 = _T_6 ? _GEN_46 : {{4'd0}, depths_13}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7798 = _T_6 ? _GEN_47 : {{4'd0}, depths_14}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7799 = _T_6 ? _GEN_48 : {{4'd0}, depths_15}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7800 = _T_6 ? _GEN_49 : {{4'd0}, depths_16}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7801 = _T_6 ? _GEN_50 : {{4'd0}, depths_17}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7802 = _T_6 ? _GEN_51 : {{4'd0}, depths_18}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7803 = _T_6 ? _GEN_52 : {{4'd0}, depths_19}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7804 = _T_6 ? _GEN_53 : {{4'd0}, depths_20}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7805 = _T_6 ? _GEN_54 : {{4'd0}, depths_21}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7806 = _T_6 ? _GEN_55 : {{4'd0}, depths_22}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7807 = _T_6 ? _GEN_56 : {{4'd0}, depths_23}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7808 = _T_6 ? _GEN_57 : {{4'd0}, depths_24}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7809 = _T_6 ? _GEN_58 : {{4'd0}, depths_25}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7810 = _T_6 ? _GEN_59 : {{4'd0}, depths_26}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7811 = _T_6 ? _GEN_60 : {{4'd0}, depths_27}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7812 = _T_6 ? _GEN_61 : {{4'd0}, depths_28}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7813 = _T_6 ? _GEN_62 : {{4'd0}, depths_29}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7814 = _T_6 ? _GEN_63 : {{4'd0}, depths_30}; // @[codewordGenerator.scala 63:27]
  wire [7:0] _GEN_7815 = _T_6 ? _GEN_64 : {{4'd0}, depths_31}; // @[codewordGenerator.scala 63:27]
  wire [30:0] _GEN_7835 = _T_6 ? {{15'd0}, _GEN_84} : _GEN_6451; // @[codewordGenerator.scala 63:27]
  assign io_outputs_codewords_0 = codewordsOut_0; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_1 = codewordsOut_1; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_2 = codewordsOut_2; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_3 = codewordsOut_3; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_4 = codewordsOut_4; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_5 = codewordsOut_5; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_6 = codewordsOut_6; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_7 = codewordsOut_7; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_8 = codewordsOut_8; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_9 = codewordsOut_9; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_10 = codewordsOut_10; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_11 = codewordsOut_11; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_12 = codewordsOut_12; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_13 = codewordsOut_13; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_14 = codewordsOut_14; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_15 = codewordsOut_15; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_16 = codewordsOut_16; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_17 = codewordsOut_17; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_18 = codewordsOut_18; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_19 = codewordsOut_19; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_20 = codewordsOut_20; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_21 = codewordsOut_21; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_22 = codewordsOut_22; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_23 = codewordsOut_23; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_24 = codewordsOut_24; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_25 = codewordsOut_25; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_26 = codewordsOut_26; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_27 = codewordsOut_27; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_28 = codewordsOut_28; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_29 = codewordsOut_29; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_30 = codewordsOut_30; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_31 = codewordsOut_31; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_32 = codewordsOut_32; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_33 = codewordsOut_33; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_34 = codewordsOut_34; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_35 = codewordsOut_35; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_36 = codewordsOut_36; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_37 = codewordsOut_37; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_38 = codewordsOut_38; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_39 = codewordsOut_39; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_40 = codewordsOut_40; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_41 = codewordsOut_41; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_42 = codewordsOut_42; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_43 = codewordsOut_43; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_44 = codewordsOut_44; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_45 = codewordsOut_45; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_46 = codewordsOut_46; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_47 = codewordsOut_47; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_48 = codewordsOut_48; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_49 = codewordsOut_49; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_50 = codewordsOut_50; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_51 = codewordsOut_51; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_52 = codewordsOut_52; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_53 = codewordsOut_53; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_54 = codewordsOut_54; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_55 = codewordsOut_55; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_56 = codewordsOut_56; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_57 = codewordsOut_57; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_58 = codewordsOut_58; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_59 = codewordsOut_59; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_60 = codewordsOut_60; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_61 = codewordsOut_61; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_62 = codewordsOut_62; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_63 = codewordsOut_63; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_64 = codewordsOut_64; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_65 = codewordsOut_65; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_66 = codewordsOut_66; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_67 = codewordsOut_67; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_68 = codewordsOut_68; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_69 = codewordsOut_69; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_70 = codewordsOut_70; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_71 = codewordsOut_71; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_72 = codewordsOut_72; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_73 = codewordsOut_73; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_74 = codewordsOut_74; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_75 = codewordsOut_75; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_76 = codewordsOut_76; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_77 = codewordsOut_77; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_78 = codewordsOut_78; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_79 = codewordsOut_79; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_80 = codewordsOut_80; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_81 = codewordsOut_81; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_82 = codewordsOut_82; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_83 = codewordsOut_83; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_84 = codewordsOut_84; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_85 = codewordsOut_85; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_86 = codewordsOut_86; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_87 = codewordsOut_87; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_88 = codewordsOut_88; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_89 = codewordsOut_89; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_90 = codewordsOut_90; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_91 = codewordsOut_91; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_92 = codewordsOut_92; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_93 = codewordsOut_93; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_94 = codewordsOut_94; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_95 = codewordsOut_95; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_96 = codewordsOut_96; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_97 = codewordsOut_97; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_98 = codewordsOut_98; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_99 = codewordsOut_99; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_100 = codewordsOut_100; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_101 = codewordsOut_101; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_102 = codewordsOut_102; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_103 = codewordsOut_103; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_104 = codewordsOut_104; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_105 = codewordsOut_105; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_106 = codewordsOut_106; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_107 = codewordsOut_107; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_108 = codewordsOut_108; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_109 = codewordsOut_109; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_110 = codewordsOut_110; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_111 = codewordsOut_111; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_112 = codewordsOut_112; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_113 = codewordsOut_113; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_114 = codewordsOut_114; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_115 = codewordsOut_115; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_116 = codewordsOut_116; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_117 = codewordsOut_117; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_118 = codewordsOut_118; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_119 = codewordsOut_119; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_120 = codewordsOut_120; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_121 = codewordsOut_121; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_122 = codewordsOut_122; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_123 = codewordsOut_123; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_124 = codewordsOut_124; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_125 = codewordsOut_125; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_126 = codewordsOut_126; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_127 = codewordsOut_127; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_128 = codewordsOut_128; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_129 = codewordsOut_129; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_130 = codewordsOut_130; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_131 = codewordsOut_131; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_132 = codewordsOut_132; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_133 = codewordsOut_133; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_134 = codewordsOut_134; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_135 = codewordsOut_135; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_136 = codewordsOut_136; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_137 = codewordsOut_137; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_138 = codewordsOut_138; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_139 = codewordsOut_139; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_140 = codewordsOut_140; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_141 = codewordsOut_141; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_142 = codewordsOut_142; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_143 = codewordsOut_143; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_144 = codewordsOut_144; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_145 = codewordsOut_145; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_146 = codewordsOut_146; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_147 = codewordsOut_147; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_148 = codewordsOut_148; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_149 = codewordsOut_149; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_150 = codewordsOut_150; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_151 = codewordsOut_151; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_152 = codewordsOut_152; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_153 = codewordsOut_153; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_154 = codewordsOut_154; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_155 = codewordsOut_155; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_156 = codewordsOut_156; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_157 = codewordsOut_157; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_158 = codewordsOut_158; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_159 = codewordsOut_159; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_160 = codewordsOut_160; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_161 = codewordsOut_161; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_162 = codewordsOut_162; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_163 = codewordsOut_163; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_164 = codewordsOut_164; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_165 = codewordsOut_165; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_166 = codewordsOut_166; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_167 = codewordsOut_167; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_168 = codewordsOut_168; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_169 = codewordsOut_169; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_170 = codewordsOut_170; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_171 = codewordsOut_171; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_172 = codewordsOut_172; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_173 = codewordsOut_173; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_174 = codewordsOut_174; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_175 = codewordsOut_175; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_176 = codewordsOut_176; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_177 = codewordsOut_177; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_178 = codewordsOut_178; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_179 = codewordsOut_179; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_180 = codewordsOut_180; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_181 = codewordsOut_181; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_182 = codewordsOut_182; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_183 = codewordsOut_183; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_184 = codewordsOut_184; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_185 = codewordsOut_185; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_186 = codewordsOut_186; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_187 = codewordsOut_187; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_188 = codewordsOut_188; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_189 = codewordsOut_189; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_190 = codewordsOut_190; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_191 = codewordsOut_191; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_192 = codewordsOut_192; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_193 = codewordsOut_193; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_194 = codewordsOut_194; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_195 = codewordsOut_195; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_196 = codewordsOut_196; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_197 = codewordsOut_197; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_198 = codewordsOut_198; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_199 = codewordsOut_199; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_200 = codewordsOut_200; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_201 = codewordsOut_201; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_202 = codewordsOut_202; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_203 = codewordsOut_203; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_204 = codewordsOut_204; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_205 = codewordsOut_205; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_206 = codewordsOut_206; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_207 = codewordsOut_207; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_208 = codewordsOut_208; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_209 = codewordsOut_209; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_210 = codewordsOut_210; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_211 = codewordsOut_211; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_212 = codewordsOut_212; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_213 = codewordsOut_213; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_214 = codewordsOut_214; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_215 = codewordsOut_215; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_216 = codewordsOut_216; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_217 = codewordsOut_217; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_218 = codewordsOut_218; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_219 = codewordsOut_219; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_220 = codewordsOut_220; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_221 = codewordsOut_221; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_222 = codewordsOut_222; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_223 = codewordsOut_223; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_224 = codewordsOut_224; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_225 = codewordsOut_225; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_226 = codewordsOut_226; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_227 = codewordsOut_227; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_228 = codewordsOut_228; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_229 = codewordsOut_229; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_230 = codewordsOut_230; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_231 = codewordsOut_231; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_232 = codewordsOut_232; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_233 = codewordsOut_233; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_234 = codewordsOut_234; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_235 = codewordsOut_235; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_236 = codewordsOut_236; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_237 = codewordsOut_237; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_238 = codewordsOut_238; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_239 = codewordsOut_239; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_240 = codewordsOut_240; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_241 = codewordsOut_241; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_242 = codewordsOut_242; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_243 = codewordsOut_243; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_244 = codewordsOut_244; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_245 = codewordsOut_245; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_246 = codewordsOut_246; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_247 = codewordsOut_247; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_248 = codewordsOut_248; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_249 = codewordsOut_249; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_250 = codewordsOut_250; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_251 = codewordsOut_251; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_252 = codewordsOut_252; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_253 = codewordsOut_253; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_254 = codewordsOut_254; // @[codewordGenerator.scala 151:24]
  assign io_outputs_codewords_255 = codewordsOut_255; // @[codewordGenerator.scala 151:24]
  assign io_outputs_lengths_0 = lengthsOut_0; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_1 = lengthsOut_1; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_2 = lengthsOut_2; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_3 = lengthsOut_3; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_4 = lengthsOut_4; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_5 = lengthsOut_5; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_6 = lengthsOut_6; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_7 = lengthsOut_7; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_8 = lengthsOut_8; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_9 = lengthsOut_9; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_10 = lengthsOut_10; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_11 = lengthsOut_11; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_12 = lengthsOut_12; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_13 = lengthsOut_13; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_14 = lengthsOut_14; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_15 = lengthsOut_15; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_16 = lengthsOut_16; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_17 = lengthsOut_17; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_18 = lengthsOut_18; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_19 = lengthsOut_19; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_20 = lengthsOut_20; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_21 = lengthsOut_21; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_22 = lengthsOut_22; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_23 = lengthsOut_23; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_24 = lengthsOut_24; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_25 = lengthsOut_25; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_26 = lengthsOut_26; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_27 = lengthsOut_27; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_28 = lengthsOut_28; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_29 = lengthsOut_29; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_30 = lengthsOut_30; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_31 = lengthsOut_31; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_32 = lengthsOut_32; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_33 = lengthsOut_33; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_34 = lengthsOut_34; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_35 = lengthsOut_35; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_36 = lengthsOut_36; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_37 = lengthsOut_37; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_38 = lengthsOut_38; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_39 = lengthsOut_39; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_40 = lengthsOut_40; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_41 = lengthsOut_41; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_42 = lengthsOut_42; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_43 = lengthsOut_43; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_44 = lengthsOut_44; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_45 = lengthsOut_45; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_46 = lengthsOut_46; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_47 = lengthsOut_47; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_48 = lengthsOut_48; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_49 = lengthsOut_49; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_50 = lengthsOut_50; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_51 = lengthsOut_51; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_52 = lengthsOut_52; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_53 = lengthsOut_53; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_54 = lengthsOut_54; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_55 = lengthsOut_55; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_56 = lengthsOut_56; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_57 = lengthsOut_57; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_58 = lengthsOut_58; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_59 = lengthsOut_59; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_60 = lengthsOut_60; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_61 = lengthsOut_61; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_62 = lengthsOut_62; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_63 = lengthsOut_63; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_64 = lengthsOut_64; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_65 = lengthsOut_65; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_66 = lengthsOut_66; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_67 = lengthsOut_67; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_68 = lengthsOut_68; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_69 = lengthsOut_69; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_70 = lengthsOut_70; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_71 = lengthsOut_71; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_72 = lengthsOut_72; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_73 = lengthsOut_73; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_74 = lengthsOut_74; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_75 = lengthsOut_75; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_76 = lengthsOut_76; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_77 = lengthsOut_77; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_78 = lengthsOut_78; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_79 = lengthsOut_79; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_80 = lengthsOut_80; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_81 = lengthsOut_81; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_82 = lengthsOut_82; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_83 = lengthsOut_83; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_84 = lengthsOut_84; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_85 = lengthsOut_85; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_86 = lengthsOut_86; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_87 = lengthsOut_87; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_88 = lengthsOut_88; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_89 = lengthsOut_89; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_90 = lengthsOut_90; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_91 = lengthsOut_91; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_92 = lengthsOut_92; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_93 = lengthsOut_93; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_94 = lengthsOut_94; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_95 = lengthsOut_95; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_96 = lengthsOut_96; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_97 = lengthsOut_97; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_98 = lengthsOut_98; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_99 = lengthsOut_99; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_100 = lengthsOut_100; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_101 = lengthsOut_101; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_102 = lengthsOut_102; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_103 = lengthsOut_103; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_104 = lengthsOut_104; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_105 = lengthsOut_105; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_106 = lengthsOut_106; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_107 = lengthsOut_107; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_108 = lengthsOut_108; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_109 = lengthsOut_109; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_110 = lengthsOut_110; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_111 = lengthsOut_111; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_112 = lengthsOut_112; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_113 = lengthsOut_113; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_114 = lengthsOut_114; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_115 = lengthsOut_115; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_116 = lengthsOut_116; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_117 = lengthsOut_117; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_118 = lengthsOut_118; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_119 = lengthsOut_119; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_120 = lengthsOut_120; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_121 = lengthsOut_121; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_122 = lengthsOut_122; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_123 = lengthsOut_123; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_124 = lengthsOut_124; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_125 = lengthsOut_125; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_126 = lengthsOut_126; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_127 = lengthsOut_127; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_128 = lengthsOut_128; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_129 = lengthsOut_129; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_130 = lengthsOut_130; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_131 = lengthsOut_131; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_132 = lengthsOut_132; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_133 = lengthsOut_133; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_134 = lengthsOut_134; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_135 = lengthsOut_135; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_136 = lengthsOut_136; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_137 = lengthsOut_137; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_138 = lengthsOut_138; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_139 = lengthsOut_139; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_140 = lengthsOut_140; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_141 = lengthsOut_141; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_142 = lengthsOut_142; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_143 = lengthsOut_143; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_144 = lengthsOut_144; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_145 = lengthsOut_145; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_146 = lengthsOut_146; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_147 = lengthsOut_147; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_148 = lengthsOut_148; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_149 = lengthsOut_149; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_150 = lengthsOut_150; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_151 = lengthsOut_151; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_152 = lengthsOut_152; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_153 = lengthsOut_153; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_154 = lengthsOut_154; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_155 = lengthsOut_155; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_156 = lengthsOut_156; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_157 = lengthsOut_157; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_158 = lengthsOut_158; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_159 = lengthsOut_159; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_160 = lengthsOut_160; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_161 = lengthsOut_161; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_162 = lengthsOut_162; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_163 = lengthsOut_163; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_164 = lengthsOut_164; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_165 = lengthsOut_165; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_166 = lengthsOut_166; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_167 = lengthsOut_167; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_168 = lengthsOut_168; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_169 = lengthsOut_169; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_170 = lengthsOut_170; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_171 = lengthsOut_171; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_172 = lengthsOut_172; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_173 = lengthsOut_173; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_174 = lengthsOut_174; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_175 = lengthsOut_175; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_176 = lengthsOut_176; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_177 = lengthsOut_177; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_178 = lengthsOut_178; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_179 = lengthsOut_179; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_180 = lengthsOut_180; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_181 = lengthsOut_181; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_182 = lengthsOut_182; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_183 = lengthsOut_183; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_184 = lengthsOut_184; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_185 = lengthsOut_185; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_186 = lengthsOut_186; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_187 = lengthsOut_187; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_188 = lengthsOut_188; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_189 = lengthsOut_189; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_190 = lengthsOut_190; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_191 = lengthsOut_191; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_192 = lengthsOut_192; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_193 = lengthsOut_193; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_194 = lengthsOut_194; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_195 = lengthsOut_195; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_196 = lengthsOut_196; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_197 = lengthsOut_197; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_198 = lengthsOut_198; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_199 = lengthsOut_199; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_200 = lengthsOut_200; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_201 = lengthsOut_201; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_202 = lengthsOut_202; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_203 = lengthsOut_203; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_204 = lengthsOut_204; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_205 = lengthsOut_205; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_206 = lengthsOut_206; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_207 = lengthsOut_207; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_208 = lengthsOut_208; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_209 = lengthsOut_209; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_210 = lengthsOut_210; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_211 = lengthsOut_211; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_212 = lengthsOut_212; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_213 = lengthsOut_213; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_214 = lengthsOut_214; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_215 = lengthsOut_215; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_216 = lengthsOut_216; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_217 = lengthsOut_217; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_218 = lengthsOut_218; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_219 = lengthsOut_219; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_220 = lengthsOut_220; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_221 = lengthsOut_221; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_222 = lengthsOut_222; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_223 = lengthsOut_223; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_224 = lengthsOut_224; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_225 = lengthsOut_225; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_226 = lengthsOut_226; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_227 = lengthsOut_227; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_228 = lengthsOut_228; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_229 = lengthsOut_229; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_230 = lengthsOut_230; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_231 = lengthsOut_231; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_232 = lengthsOut_232; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_233 = lengthsOut_233; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_234 = lengthsOut_234; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_235 = lengthsOut_235; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_236 = lengthsOut_236; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_237 = lengthsOut_237; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_238 = lengthsOut_238; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_239 = lengthsOut_239; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_240 = lengthsOut_240; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_241 = lengthsOut_241; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_242 = lengthsOut_242; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_243 = lengthsOut_243; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_244 = lengthsOut_244; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_245 = lengthsOut_245; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_246 = lengthsOut_246; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_247 = lengthsOut_247; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_248 = lengthsOut_248; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_249 = lengthsOut_249; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_250 = lengthsOut_250; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_251 = lengthsOut_251; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_252 = lengthsOut_252; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_253 = lengthsOut_253; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_254 = lengthsOut_254; // @[codewordGenerator.scala 152:22]
  assign io_outputs_lengths_255 = lengthsOut_255; // @[codewordGenerator.scala 152:22]
  assign io_outputs_charactersOut_0 = charactersIn_0; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_1 = charactersIn_1; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_2 = charactersIn_2; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_3 = charactersIn_3; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_4 = charactersIn_4; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_5 = charactersIn_5; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_6 = charactersIn_6; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_7 = charactersIn_7; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_8 = charactersIn_8; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_9 = charactersIn_9; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_10 = charactersIn_10; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_11 = charactersIn_11; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_12 = charactersIn_12; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_13 = charactersIn_13; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_14 = charactersIn_14; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_15 = charactersIn_15; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_16 = charactersIn_16; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_17 = charactersIn_17; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_18 = charactersIn_18; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_19 = charactersIn_19; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_20 = charactersIn_20; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_21 = charactersIn_21; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_22 = charactersIn_22; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_23 = charactersIn_23; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_24 = charactersIn_24; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_25 = charactersIn_25; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_26 = charactersIn_26; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_27 = charactersIn_27; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_28 = charactersIn_28; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_29 = charactersIn_29; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_30 = charactersIn_30; // @[codewordGenerator.scala 153:28]
  assign io_outputs_charactersOut_31 = charactersIn_31; // @[codewordGenerator.scala 153:28]
  assign io_outputs_nodes = nodes; // @[codewordGenerator.scala 154:20]
  assign io_outputs_escapeCharacterLength = escapeCharacterLength; // @[codewordGenerator.scala 156:36]
  assign io_outputs_escapeCodeword = escapeCodeword; // @[codewordGenerator.scala 159:29]
  assign io_finished = state == 2'h0; // @[codewordGenerator.scala 160:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  charactersIn_0 = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  charactersIn_1 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  charactersIn_2 = _RAND_3[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  charactersIn_3 = _RAND_4[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  charactersIn_4 = _RAND_5[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  charactersIn_5 = _RAND_6[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  charactersIn_6 = _RAND_7[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  charactersIn_7 = _RAND_8[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  charactersIn_8 = _RAND_9[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  charactersIn_9 = _RAND_10[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  charactersIn_10 = _RAND_11[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  charactersIn_11 = _RAND_12[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  charactersIn_12 = _RAND_13[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  charactersIn_13 = _RAND_14[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  charactersIn_14 = _RAND_15[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  charactersIn_15 = _RAND_16[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  charactersIn_16 = _RAND_17[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  charactersIn_17 = _RAND_18[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  charactersIn_18 = _RAND_19[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  charactersIn_19 = _RAND_20[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  charactersIn_20 = _RAND_21[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  charactersIn_21 = _RAND_22[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  charactersIn_22 = _RAND_23[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  charactersIn_23 = _RAND_24[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  charactersIn_24 = _RAND_25[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  charactersIn_25 = _RAND_26[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  charactersIn_26 = _RAND_27[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  charactersIn_27 = _RAND_28[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  charactersIn_28 = _RAND_29[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  charactersIn_29 = _RAND_30[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  charactersIn_30 = _RAND_31[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  charactersIn_31 = _RAND_32[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  depths_0 = _RAND_33[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  depths_1 = _RAND_34[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  depths_2 = _RAND_35[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  depths_3 = _RAND_36[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  depths_4 = _RAND_37[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  depths_5 = _RAND_38[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  depths_6 = _RAND_39[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  depths_7 = _RAND_40[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  depths_8 = _RAND_41[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  depths_9 = _RAND_42[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  depths_10 = _RAND_43[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  depths_11 = _RAND_44[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  depths_12 = _RAND_45[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  depths_13 = _RAND_46[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  depths_14 = _RAND_47[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  depths_15 = _RAND_48[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  depths_16 = _RAND_49[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  depths_17 = _RAND_50[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  depths_18 = _RAND_51[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  depths_19 = _RAND_52[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  depths_20 = _RAND_53[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  depths_21 = _RAND_54[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  depths_22 = _RAND_55[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  depths_23 = _RAND_56[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  depths_24 = _RAND_57[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  depths_25 = _RAND_58[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  depths_26 = _RAND_59[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  depths_27 = _RAND_60[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  depths_28 = _RAND_61[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  depths_29 = _RAND_62[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  depths_30 = _RAND_63[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  depths_31 = _RAND_64[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  codewords_0 = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  codewords_1 = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  codewords_2 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  codewords_3 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  codewords_4 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  codewords_5 = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  codewords_6 = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  codewords_7 = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  codewords_8 = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  codewords_9 = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  codewords_10 = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  codewords_11 = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  codewords_12 = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  codewords_13 = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  codewords_14 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  codewords_15 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  codewords_16 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  codewords_17 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  codewords_18 = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  codewords_19 = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  codewords_20 = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  codewords_21 = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  codewords_22 = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  codewords_23 = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  codewords_24 = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  codewords_25 = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  codewords_26 = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  codewords_27 = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  codewords_28 = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  codewords_29 = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  codewords_30 = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  codewords_31 = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  codewords_32 = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  codewords_33 = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  codewords_34 = _RAND_99[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  codewords_35 = _RAND_100[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  codewords_36 = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  codewords_37 = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  codewords_38 = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  codewords_39 = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  codewords_40 = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  codewords_41 = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  codewords_42 = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  codewords_43 = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  codewords_44 = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  codewords_45 = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  codewords_46 = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  codewords_47 = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  codewords_48 = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  codewords_49 = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  codewords_50 = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  codewords_51 = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  codewords_52 = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  codewords_53 = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  codewords_54 = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  codewords_55 = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  codewords_56 = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  codewords_57 = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  codewords_58 = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  codewords_59 = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  codewords_60 = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  codewords_61 = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  codewords_62 = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  codewords_63 = _RAND_128[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  codewords_64 = _RAND_129[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  codewords_65 = _RAND_130[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  codewords_66 = _RAND_131[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  codewords_67 = _RAND_132[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  codewords_68 = _RAND_133[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  codewords_69 = _RAND_134[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  codewords_70 = _RAND_135[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  codewords_71 = _RAND_136[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  codewords_72 = _RAND_137[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  codewords_73 = _RAND_138[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  codewords_74 = _RAND_139[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  codewords_75 = _RAND_140[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  codewords_76 = _RAND_141[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  codewords_77 = _RAND_142[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  codewords_78 = _RAND_143[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  codewords_79 = _RAND_144[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  codewords_80 = _RAND_145[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  codewords_81 = _RAND_146[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  codewords_82 = _RAND_147[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  codewords_83 = _RAND_148[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  codewords_84 = _RAND_149[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  codewords_85 = _RAND_150[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  codewords_86 = _RAND_151[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  codewords_87 = _RAND_152[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  codewords_88 = _RAND_153[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  codewords_89 = _RAND_154[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  codewords_90 = _RAND_155[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  codewords_91 = _RAND_156[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  codewords_92 = _RAND_157[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  codewords_93 = _RAND_158[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  codewords_94 = _RAND_159[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  codewords_95 = _RAND_160[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  codewords_96 = _RAND_161[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  codewords_97 = _RAND_162[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  codewords_98 = _RAND_163[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  codewords_99 = _RAND_164[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  codewords_100 = _RAND_165[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  codewords_101 = _RAND_166[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  codewords_102 = _RAND_167[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  codewords_103 = _RAND_168[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  codewords_104 = _RAND_169[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  codewords_105 = _RAND_170[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  codewords_106 = _RAND_171[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  codewords_107 = _RAND_172[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  codewords_108 = _RAND_173[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  codewords_109 = _RAND_174[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  codewords_110 = _RAND_175[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  codewords_111 = _RAND_176[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  codewords_112 = _RAND_177[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  codewords_113 = _RAND_178[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  codewords_114 = _RAND_179[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  codewords_115 = _RAND_180[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  codewords_116 = _RAND_181[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  codewords_117 = _RAND_182[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  codewords_118 = _RAND_183[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  codewords_119 = _RAND_184[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  codewords_120 = _RAND_185[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  codewords_121 = _RAND_186[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  codewords_122 = _RAND_187[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  codewords_123 = _RAND_188[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  codewords_124 = _RAND_189[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  codewords_125 = _RAND_190[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  codewords_126 = _RAND_191[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  codewords_127 = _RAND_192[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  codewords_128 = _RAND_193[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  codewords_129 = _RAND_194[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  codewords_130 = _RAND_195[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  codewords_131 = _RAND_196[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  codewords_132 = _RAND_197[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  codewords_133 = _RAND_198[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  codewords_134 = _RAND_199[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  codewords_135 = _RAND_200[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  codewords_136 = _RAND_201[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  codewords_137 = _RAND_202[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  codewords_138 = _RAND_203[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  codewords_139 = _RAND_204[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  codewords_140 = _RAND_205[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  codewords_141 = _RAND_206[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  codewords_142 = _RAND_207[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  codewords_143 = _RAND_208[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  codewords_144 = _RAND_209[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  codewords_145 = _RAND_210[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  codewords_146 = _RAND_211[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  codewords_147 = _RAND_212[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  codewords_148 = _RAND_213[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  codewords_149 = _RAND_214[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  codewords_150 = _RAND_215[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  codewords_151 = _RAND_216[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  codewords_152 = _RAND_217[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  codewords_153 = _RAND_218[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  codewords_154 = _RAND_219[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  codewords_155 = _RAND_220[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  codewords_156 = _RAND_221[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  codewords_157 = _RAND_222[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  codewords_158 = _RAND_223[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  codewords_159 = _RAND_224[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  codewords_160 = _RAND_225[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  codewords_161 = _RAND_226[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  codewords_162 = _RAND_227[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  codewords_163 = _RAND_228[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  codewords_164 = _RAND_229[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  codewords_165 = _RAND_230[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  codewords_166 = _RAND_231[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  codewords_167 = _RAND_232[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  codewords_168 = _RAND_233[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  codewords_169 = _RAND_234[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  codewords_170 = _RAND_235[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  codewords_171 = _RAND_236[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  codewords_172 = _RAND_237[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  codewords_173 = _RAND_238[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  codewords_174 = _RAND_239[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  codewords_175 = _RAND_240[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  codewords_176 = _RAND_241[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  codewords_177 = _RAND_242[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  codewords_178 = _RAND_243[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  codewords_179 = _RAND_244[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  codewords_180 = _RAND_245[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  codewords_181 = _RAND_246[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  codewords_182 = _RAND_247[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  codewords_183 = _RAND_248[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  codewords_184 = _RAND_249[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  codewords_185 = _RAND_250[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  codewords_186 = _RAND_251[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  codewords_187 = _RAND_252[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  codewords_188 = _RAND_253[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  codewords_189 = _RAND_254[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  codewords_190 = _RAND_255[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  codewords_191 = _RAND_256[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  codewords_192 = _RAND_257[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  codewords_193 = _RAND_258[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  codewords_194 = _RAND_259[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  codewords_195 = _RAND_260[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  codewords_196 = _RAND_261[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  codewords_197 = _RAND_262[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  codewords_198 = _RAND_263[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  codewords_199 = _RAND_264[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  codewords_200 = _RAND_265[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  codewords_201 = _RAND_266[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  codewords_202 = _RAND_267[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  codewords_203 = _RAND_268[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  codewords_204 = _RAND_269[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  codewords_205 = _RAND_270[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  codewords_206 = _RAND_271[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  codewords_207 = _RAND_272[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  codewords_208 = _RAND_273[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  codewords_209 = _RAND_274[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  codewords_210 = _RAND_275[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  codewords_211 = _RAND_276[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  codewords_212 = _RAND_277[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  codewords_213 = _RAND_278[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  codewords_214 = _RAND_279[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  codewords_215 = _RAND_280[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  codewords_216 = _RAND_281[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  codewords_217 = _RAND_282[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  codewords_218 = _RAND_283[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  codewords_219 = _RAND_284[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  codewords_220 = _RAND_285[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  codewords_221 = _RAND_286[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  codewords_222 = _RAND_287[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  codewords_223 = _RAND_288[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  codewords_224 = _RAND_289[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  codewords_225 = _RAND_290[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  codewords_226 = _RAND_291[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  codewords_227 = _RAND_292[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  codewords_228 = _RAND_293[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  codewords_229 = _RAND_294[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  codewords_230 = _RAND_295[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  codewords_231 = _RAND_296[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  codewords_232 = _RAND_297[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  codewords_233 = _RAND_298[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  codewords_234 = _RAND_299[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  codewords_235 = _RAND_300[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  codewords_236 = _RAND_301[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  codewords_237 = _RAND_302[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  codewords_238 = _RAND_303[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  codewords_239 = _RAND_304[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  codewords_240 = _RAND_305[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  codewords_241 = _RAND_306[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  codewords_242 = _RAND_307[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  codewords_243 = _RAND_308[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  codewords_244 = _RAND_309[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  codewords_245 = _RAND_310[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  codewords_246 = _RAND_311[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  codewords_247 = _RAND_312[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  codewords_248 = _RAND_313[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  codewords_249 = _RAND_314[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  codewords_250 = _RAND_315[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  codewords_251 = _RAND_316[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  codewords_252 = _RAND_317[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  codewords_253 = _RAND_318[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  codewords_254 = _RAND_319[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  codewords_255 = _RAND_320[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  codewordsOut_0 = _RAND_321[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  codewordsOut_1 = _RAND_322[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  codewordsOut_2 = _RAND_323[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  codewordsOut_3 = _RAND_324[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  codewordsOut_4 = _RAND_325[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  codewordsOut_5 = _RAND_326[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  codewordsOut_6 = _RAND_327[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  codewordsOut_7 = _RAND_328[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  codewordsOut_8 = _RAND_329[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  codewordsOut_9 = _RAND_330[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  codewordsOut_10 = _RAND_331[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  codewordsOut_11 = _RAND_332[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  codewordsOut_12 = _RAND_333[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  codewordsOut_13 = _RAND_334[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  codewordsOut_14 = _RAND_335[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  codewordsOut_15 = _RAND_336[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  codewordsOut_16 = _RAND_337[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  codewordsOut_17 = _RAND_338[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  codewordsOut_18 = _RAND_339[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  codewordsOut_19 = _RAND_340[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  codewordsOut_20 = _RAND_341[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  codewordsOut_21 = _RAND_342[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  codewordsOut_22 = _RAND_343[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  codewordsOut_23 = _RAND_344[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  codewordsOut_24 = _RAND_345[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  codewordsOut_25 = _RAND_346[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  codewordsOut_26 = _RAND_347[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  codewordsOut_27 = _RAND_348[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  codewordsOut_28 = _RAND_349[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  codewordsOut_29 = _RAND_350[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  codewordsOut_30 = _RAND_351[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  codewordsOut_31 = _RAND_352[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  codewordsOut_32 = _RAND_353[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  codewordsOut_33 = _RAND_354[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  codewordsOut_34 = _RAND_355[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  codewordsOut_35 = _RAND_356[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  codewordsOut_36 = _RAND_357[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  codewordsOut_37 = _RAND_358[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  codewordsOut_38 = _RAND_359[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  codewordsOut_39 = _RAND_360[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  codewordsOut_40 = _RAND_361[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  codewordsOut_41 = _RAND_362[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  codewordsOut_42 = _RAND_363[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  codewordsOut_43 = _RAND_364[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  codewordsOut_44 = _RAND_365[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  codewordsOut_45 = _RAND_366[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  codewordsOut_46 = _RAND_367[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  codewordsOut_47 = _RAND_368[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  codewordsOut_48 = _RAND_369[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  codewordsOut_49 = _RAND_370[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  codewordsOut_50 = _RAND_371[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  codewordsOut_51 = _RAND_372[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  codewordsOut_52 = _RAND_373[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  codewordsOut_53 = _RAND_374[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  codewordsOut_54 = _RAND_375[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  codewordsOut_55 = _RAND_376[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  codewordsOut_56 = _RAND_377[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  codewordsOut_57 = _RAND_378[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  codewordsOut_58 = _RAND_379[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  codewordsOut_59 = _RAND_380[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  codewordsOut_60 = _RAND_381[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  codewordsOut_61 = _RAND_382[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  codewordsOut_62 = _RAND_383[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  codewordsOut_63 = _RAND_384[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  codewordsOut_64 = _RAND_385[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  codewordsOut_65 = _RAND_386[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  codewordsOut_66 = _RAND_387[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  codewordsOut_67 = _RAND_388[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  codewordsOut_68 = _RAND_389[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  codewordsOut_69 = _RAND_390[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  codewordsOut_70 = _RAND_391[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  codewordsOut_71 = _RAND_392[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  codewordsOut_72 = _RAND_393[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  codewordsOut_73 = _RAND_394[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  codewordsOut_74 = _RAND_395[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  codewordsOut_75 = _RAND_396[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  codewordsOut_76 = _RAND_397[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  codewordsOut_77 = _RAND_398[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  codewordsOut_78 = _RAND_399[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  codewordsOut_79 = _RAND_400[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  codewordsOut_80 = _RAND_401[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  codewordsOut_81 = _RAND_402[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  codewordsOut_82 = _RAND_403[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  codewordsOut_83 = _RAND_404[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  codewordsOut_84 = _RAND_405[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  codewordsOut_85 = _RAND_406[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  codewordsOut_86 = _RAND_407[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  codewordsOut_87 = _RAND_408[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  codewordsOut_88 = _RAND_409[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  codewordsOut_89 = _RAND_410[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  codewordsOut_90 = _RAND_411[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  codewordsOut_91 = _RAND_412[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  codewordsOut_92 = _RAND_413[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  codewordsOut_93 = _RAND_414[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  codewordsOut_94 = _RAND_415[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  codewordsOut_95 = _RAND_416[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  codewordsOut_96 = _RAND_417[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  codewordsOut_97 = _RAND_418[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  codewordsOut_98 = _RAND_419[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  codewordsOut_99 = _RAND_420[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  codewordsOut_100 = _RAND_421[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  codewordsOut_101 = _RAND_422[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  codewordsOut_102 = _RAND_423[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  codewordsOut_103 = _RAND_424[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  codewordsOut_104 = _RAND_425[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  codewordsOut_105 = _RAND_426[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  codewordsOut_106 = _RAND_427[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  codewordsOut_107 = _RAND_428[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  codewordsOut_108 = _RAND_429[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  codewordsOut_109 = _RAND_430[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  codewordsOut_110 = _RAND_431[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  codewordsOut_111 = _RAND_432[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  codewordsOut_112 = _RAND_433[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  codewordsOut_113 = _RAND_434[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  codewordsOut_114 = _RAND_435[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  codewordsOut_115 = _RAND_436[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  codewordsOut_116 = _RAND_437[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  codewordsOut_117 = _RAND_438[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  codewordsOut_118 = _RAND_439[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  codewordsOut_119 = _RAND_440[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  codewordsOut_120 = _RAND_441[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  codewordsOut_121 = _RAND_442[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  codewordsOut_122 = _RAND_443[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  codewordsOut_123 = _RAND_444[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  codewordsOut_124 = _RAND_445[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  codewordsOut_125 = _RAND_446[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  codewordsOut_126 = _RAND_447[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  codewordsOut_127 = _RAND_448[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  codewordsOut_128 = _RAND_449[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  codewordsOut_129 = _RAND_450[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  codewordsOut_130 = _RAND_451[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  codewordsOut_131 = _RAND_452[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  codewordsOut_132 = _RAND_453[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  codewordsOut_133 = _RAND_454[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  codewordsOut_134 = _RAND_455[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  codewordsOut_135 = _RAND_456[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  codewordsOut_136 = _RAND_457[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  codewordsOut_137 = _RAND_458[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  codewordsOut_138 = _RAND_459[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  codewordsOut_139 = _RAND_460[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  codewordsOut_140 = _RAND_461[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  codewordsOut_141 = _RAND_462[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  codewordsOut_142 = _RAND_463[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  codewordsOut_143 = _RAND_464[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  codewordsOut_144 = _RAND_465[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  codewordsOut_145 = _RAND_466[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  codewordsOut_146 = _RAND_467[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  codewordsOut_147 = _RAND_468[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  codewordsOut_148 = _RAND_469[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  codewordsOut_149 = _RAND_470[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  codewordsOut_150 = _RAND_471[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  codewordsOut_151 = _RAND_472[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  codewordsOut_152 = _RAND_473[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  codewordsOut_153 = _RAND_474[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  codewordsOut_154 = _RAND_475[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  codewordsOut_155 = _RAND_476[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  codewordsOut_156 = _RAND_477[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  codewordsOut_157 = _RAND_478[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  codewordsOut_158 = _RAND_479[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  codewordsOut_159 = _RAND_480[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  codewordsOut_160 = _RAND_481[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  codewordsOut_161 = _RAND_482[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  codewordsOut_162 = _RAND_483[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  codewordsOut_163 = _RAND_484[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  codewordsOut_164 = _RAND_485[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  codewordsOut_165 = _RAND_486[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  codewordsOut_166 = _RAND_487[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  codewordsOut_167 = _RAND_488[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  codewordsOut_168 = _RAND_489[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  codewordsOut_169 = _RAND_490[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  codewordsOut_170 = _RAND_491[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  codewordsOut_171 = _RAND_492[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  codewordsOut_172 = _RAND_493[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  codewordsOut_173 = _RAND_494[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  codewordsOut_174 = _RAND_495[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  codewordsOut_175 = _RAND_496[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  codewordsOut_176 = _RAND_497[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  codewordsOut_177 = _RAND_498[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  codewordsOut_178 = _RAND_499[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  codewordsOut_179 = _RAND_500[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  codewordsOut_180 = _RAND_501[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  codewordsOut_181 = _RAND_502[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  codewordsOut_182 = _RAND_503[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  codewordsOut_183 = _RAND_504[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  codewordsOut_184 = _RAND_505[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  codewordsOut_185 = _RAND_506[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  codewordsOut_186 = _RAND_507[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  codewordsOut_187 = _RAND_508[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  codewordsOut_188 = _RAND_509[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  codewordsOut_189 = _RAND_510[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  codewordsOut_190 = _RAND_511[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  codewordsOut_191 = _RAND_512[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  codewordsOut_192 = _RAND_513[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  codewordsOut_193 = _RAND_514[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  codewordsOut_194 = _RAND_515[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  codewordsOut_195 = _RAND_516[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  codewordsOut_196 = _RAND_517[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  codewordsOut_197 = _RAND_518[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  codewordsOut_198 = _RAND_519[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  codewordsOut_199 = _RAND_520[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  codewordsOut_200 = _RAND_521[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  codewordsOut_201 = _RAND_522[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  codewordsOut_202 = _RAND_523[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  codewordsOut_203 = _RAND_524[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  codewordsOut_204 = _RAND_525[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  codewordsOut_205 = _RAND_526[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  codewordsOut_206 = _RAND_527[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  codewordsOut_207 = _RAND_528[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  codewordsOut_208 = _RAND_529[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  codewordsOut_209 = _RAND_530[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  codewordsOut_210 = _RAND_531[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  codewordsOut_211 = _RAND_532[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  codewordsOut_212 = _RAND_533[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  codewordsOut_213 = _RAND_534[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  codewordsOut_214 = _RAND_535[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  codewordsOut_215 = _RAND_536[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  codewordsOut_216 = _RAND_537[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  codewordsOut_217 = _RAND_538[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  codewordsOut_218 = _RAND_539[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  codewordsOut_219 = _RAND_540[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  codewordsOut_220 = _RAND_541[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  codewordsOut_221 = _RAND_542[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  codewordsOut_222 = _RAND_543[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  codewordsOut_223 = _RAND_544[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  codewordsOut_224 = _RAND_545[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  codewordsOut_225 = _RAND_546[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  codewordsOut_226 = _RAND_547[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  codewordsOut_227 = _RAND_548[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  codewordsOut_228 = _RAND_549[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  codewordsOut_229 = _RAND_550[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  codewordsOut_230 = _RAND_551[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  codewordsOut_231 = _RAND_552[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  codewordsOut_232 = _RAND_553[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  codewordsOut_233 = _RAND_554[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  codewordsOut_234 = _RAND_555[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  codewordsOut_235 = _RAND_556[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  codewordsOut_236 = _RAND_557[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  codewordsOut_237 = _RAND_558[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  codewordsOut_238 = _RAND_559[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  codewordsOut_239 = _RAND_560[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  codewordsOut_240 = _RAND_561[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  codewordsOut_241 = _RAND_562[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  codewordsOut_242 = _RAND_563[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  codewordsOut_243 = _RAND_564[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  codewordsOut_244 = _RAND_565[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  codewordsOut_245 = _RAND_566[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  codewordsOut_246 = _RAND_567[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  codewordsOut_247 = _RAND_568[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  codewordsOut_248 = _RAND_569[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  codewordsOut_249 = _RAND_570[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  codewordsOut_250 = _RAND_571[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  codewordsOut_251 = _RAND_572[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  codewordsOut_252 = _RAND_573[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  codewordsOut_253 = _RAND_574[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  codewordsOut_254 = _RAND_575[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  codewordsOut_255 = _RAND_576[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  lengths_0 = _RAND_577[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  lengths_1 = _RAND_578[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  lengths_2 = _RAND_579[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  lengths_3 = _RAND_580[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  lengths_4 = _RAND_581[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  lengths_5 = _RAND_582[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  lengths_6 = _RAND_583[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  lengths_7 = _RAND_584[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  lengths_8 = _RAND_585[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  lengths_9 = _RAND_586[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  lengths_10 = _RAND_587[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  lengths_11 = _RAND_588[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  lengths_12 = _RAND_589[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  lengths_13 = _RAND_590[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  lengths_14 = _RAND_591[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  lengths_15 = _RAND_592[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  lengths_16 = _RAND_593[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  lengths_17 = _RAND_594[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  lengths_18 = _RAND_595[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  lengths_19 = _RAND_596[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  lengths_20 = _RAND_597[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  lengths_21 = _RAND_598[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  lengths_22 = _RAND_599[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  lengths_23 = _RAND_600[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  lengths_24 = _RAND_601[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  lengths_25 = _RAND_602[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  lengths_26 = _RAND_603[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  lengths_27 = _RAND_604[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  lengths_28 = _RAND_605[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  lengths_29 = _RAND_606[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  lengths_30 = _RAND_607[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  lengths_31 = _RAND_608[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  lengths_32 = _RAND_609[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  lengths_33 = _RAND_610[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  lengths_34 = _RAND_611[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  lengths_35 = _RAND_612[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  lengths_36 = _RAND_613[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  lengths_37 = _RAND_614[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  lengths_38 = _RAND_615[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  lengths_39 = _RAND_616[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  lengths_40 = _RAND_617[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  lengths_41 = _RAND_618[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  lengths_42 = _RAND_619[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  lengths_43 = _RAND_620[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  lengths_44 = _RAND_621[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  lengths_45 = _RAND_622[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  lengths_46 = _RAND_623[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  lengths_47 = _RAND_624[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  lengths_48 = _RAND_625[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  lengths_49 = _RAND_626[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  lengths_50 = _RAND_627[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  lengths_51 = _RAND_628[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  lengths_52 = _RAND_629[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  lengths_53 = _RAND_630[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  lengths_54 = _RAND_631[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  lengths_55 = _RAND_632[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  lengths_56 = _RAND_633[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  lengths_57 = _RAND_634[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  lengths_58 = _RAND_635[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  lengths_59 = _RAND_636[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  lengths_60 = _RAND_637[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  lengths_61 = _RAND_638[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  lengths_62 = _RAND_639[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  lengths_63 = _RAND_640[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  lengths_64 = _RAND_641[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  lengths_65 = _RAND_642[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  lengths_66 = _RAND_643[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  lengths_67 = _RAND_644[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  lengths_68 = _RAND_645[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  lengths_69 = _RAND_646[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  lengths_70 = _RAND_647[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  lengths_71 = _RAND_648[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  lengths_72 = _RAND_649[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  lengths_73 = _RAND_650[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  lengths_74 = _RAND_651[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  lengths_75 = _RAND_652[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  lengths_76 = _RAND_653[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  lengths_77 = _RAND_654[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  lengths_78 = _RAND_655[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  lengths_79 = _RAND_656[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  lengths_80 = _RAND_657[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  lengths_81 = _RAND_658[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  lengths_82 = _RAND_659[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  lengths_83 = _RAND_660[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  lengths_84 = _RAND_661[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  lengths_85 = _RAND_662[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  lengths_86 = _RAND_663[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  lengths_87 = _RAND_664[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  lengths_88 = _RAND_665[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  lengths_89 = _RAND_666[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  lengths_90 = _RAND_667[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  lengths_91 = _RAND_668[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  lengths_92 = _RAND_669[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  lengths_93 = _RAND_670[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  lengths_94 = _RAND_671[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  lengths_95 = _RAND_672[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  lengths_96 = _RAND_673[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  lengths_97 = _RAND_674[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  lengths_98 = _RAND_675[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  lengths_99 = _RAND_676[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  lengths_100 = _RAND_677[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  lengths_101 = _RAND_678[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  lengths_102 = _RAND_679[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  lengths_103 = _RAND_680[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  lengths_104 = _RAND_681[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{`RANDOM}};
  lengths_105 = _RAND_682[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  lengths_106 = _RAND_683[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  lengths_107 = _RAND_684[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  lengths_108 = _RAND_685[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  lengths_109 = _RAND_686[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  lengths_110 = _RAND_687[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  lengths_111 = _RAND_688[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  lengths_112 = _RAND_689[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  lengths_113 = _RAND_690[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  lengths_114 = _RAND_691[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  lengths_115 = _RAND_692[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  lengths_116 = _RAND_693[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  lengths_117 = _RAND_694[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  lengths_118 = _RAND_695[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  lengths_119 = _RAND_696[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  lengths_120 = _RAND_697[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  lengths_121 = _RAND_698[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  lengths_122 = _RAND_699[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  lengths_123 = _RAND_700[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  lengths_124 = _RAND_701[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  lengths_125 = _RAND_702[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  lengths_126 = _RAND_703[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  lengths_127 = _RAND_704[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  lengths_128 = _RAND_705[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  lengths_129 = _RAND_706[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  lengths_130 = _RAND_707[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  lengths_131 = _RAND_708[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  lengths_132 = _RAND_709[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  lengths_133 = _RAND_710[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  lengths_134 = _RAND_711[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  lengths_135 = _RAND_712[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  lengths_136 = _RAND_713[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  lengths_137 = _RAND_714[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  lengths_138 = _RAND_715[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  lengths_139 = _RAND_716[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  lengths_140 = _RAND_717[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  lengths_141 = _RAND_718[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  lengths_142 = _RAND_719[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  lengths_143 = _RAND_720[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  lengths_144 = _RAND_721[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  lengths_145 = _RAND_722[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{`RANDOM}};
  lengths_146 = _RAND_723[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{`RANDOM}};
  lengths_147 = _RAND_724[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{`RANDOM}};
  lengths_148 = _RAND_725[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{`RANDOM}};
  lengths_149 = _RAND_726[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{`RANDOM}};
  lengths_150 = _RAND_727[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{`RANDOM}};
  lengths_151 = _RAND_728[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{`RANDOM}};
  lengths_152 = _RAND_729[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{`RANDOM}};
  lengths_153 = _RAND_730[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{`RANDOM}};
  lengths_154 = _RAND_731[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{`RANDOM}};
  lengths_155 = _RAND_732[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{`RANDOM}};
  lengths_156 = _RAND_733[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{`RANDOM}};
  lengths_157 = _RAND_734[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{`RANDOM}};
  lengths_158 = _RAND_735[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{`RANDOM}};
  lengths_159 = _RAND_736[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{`RANDOM}};
  lengths_160 = _RAND_737[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{`RANDOM}};
  lengths_161 = _RAND_738[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{`RANDOM}};
  lengths_162 = _RAND_739[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{`RANDOM}};
  lengths_163 = _RAND_740[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{`RANDOM}};
  lengths_164 = _RAND_741[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{`RANDOM}};
  lengths_165 = _RAND_742[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{`RANDOM}};
  lengths_166 = _RAND_743[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{`RANDOM}};
  lengths_167 = _RAND_744[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{`RANDOM}};
  lengths_168 = _RAND_745[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{`RANDOM}};
  lengths_169 = _RAND_746[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{`RANDOM}};
  lengths_170 = _RAND_747[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{`RANDOM}};
  lengths_171 = _RAND_748[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{`RANDOM}};
  lengths_172 = _RAND_749[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{`RANDOM}};
  lengths_173 = _RAND_750[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{`RANDOM}};
  lengths_174 = _RAND_751[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{`RANDOM}};
  lengths_175 = _RAND_752[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{`RANDOM}};
  lengths_176 = _RAND_753[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{`RANDOM}};
  lengths_177 = _RAND_754[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_755 = {1{`RANDOM}};
  lengths_178 = _RAND_755[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_756 = {1{`RANDOM}};
  lengths_179 = _RAND_756[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_757 = {1{`RANDOM}};
  lengths_180 = _RAND_757[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_758 = {1{`RANDOM}};
  lengths_181 = _RAND_758[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_759 = {1{`RANDOM}};
  lengths_182 = _RAND_759[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_760 = {1{`RANDOM}};
  lengths_183 = _RAND_760[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_761 = {1{`RANDOM}};
  lengths_184 = _RAND_761[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_762 = {1{`RANDOM}};
  lengths_185 = _RAND_762[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_763 = {1{`RANDOM}};
  lengths_186 = _RAND_763[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_764 = {1{`RANDOM}};
  lengths_187 = _RAND_764[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_765 = {1{`RANDOM}};
  lengths_188 = _RAND_765[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_766 = {1{`RANDOM}};
  lengths_189 = _RAND_766[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_767 = {1{`RANDOM}};
  lengths_190 = _RAND_767[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_768 = {1{`RANDOM}};
  lengths_191 = _RAND_768[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_769 = {1{`RANDOM}};
  lengths_192 = _RAND_769[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_770 = {1{`RANDOM}};
  lengths_193 = _RAND_770[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_771 = {1{`RANDOM}};
  lengths_194 = _RAND_771[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_772 = {1{`RANDOM}};
  lengths_195 = _RAND_772[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_773 = {1{`RANDOM}};
  lengths_196 = _RAND_773[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_774 = {1{`RANDOM}};
  lengths_197 = _RAND_774[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_775 = {1{`RANDOM}};
  lengths_198 = _RAND_775[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_776 = {1{`RANDOM}};
  lengths_199 = _RAND_776[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_777 = {1{`RANDOM}};
  lengths_200 = _RAND_777[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_778 = {1{`RANDOM}};
  lengths_201 = _RAND_778[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_779 = {1{`RANDOM}};
  lengths_202 = _RAND_779[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_780 = {1{`RANDOM}};
  lengths_203 = _RAND_780[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_781 = {1{`RANDOM}};
  lengths_204 = _RAND_781[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_782 = {1{`RANDOM}};
  lengths_205 = _RAND_782[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_783 = {1{`RANDOM}};
  lengths_206 = _RAND_783[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_784 = {1{`RANDOM}};
  lengths_207 = _RAND_784[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_785 = {1{`RANDOM}};
  lengths_208 = _RAND_785[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_786 = {1{`RANDOM}};
  lengths_209 = _RAND_786[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_787 = {1{`RANDOM}};
  lengths_210 = _RAND_787[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_788 = {1{`RANDOM}};
  lengths_211 = _RAND_788[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_789 = {1{`RANDOM}};
  lengths_212 = _RAND_789[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_790 = {1{`RANDOM}};
  lengths_213 = _RAND_790[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_791 = {1{`RANDOM}};
  lengths_214 = _RAND_791[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_792 = {1{`RANDOM}};
  lengths_215 = _RAND_792[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_793 = {1{`RANDOM}};
  lengths_216 = _RAND_793[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_794 = {1{`RANDOM}};
  lengths_217 = _RAND_794[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_795 = {1{`RANDOM}};
  lengths_218 = _RAND_795[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_796 = {1{`RANDOM}};
  lengths_219 = _RAND_796[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_797 = {1{`RANDOM}};
  lengths_220 = _RAND_797[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_798 = {1{`RANDOM}};
  lengths_221 = _RAND_798[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_799 = {1{`RANDOM}};
  lengths_222 = _RAND_799[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_800 = {1{`RANDOM}};
  lengths_223 = _RAND_800[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_801 = {1{`RANDOM}};
  lengths_224 = _RAND_801[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_802 = {1{`RANDOM}};
  lengths_225 = _RAND_802[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_803 = {1{`RANDOM}};
  lengths_226 = _RAND_803[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_804 = {1{`RANDOM}};
  lengths_227 = _RAND_804[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_805 = {1{`RANDOM}};
  lengths_228 = _RAND_805[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_806 = {1{`RANDOM}};
  lengths_229 = _RAND_806[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_807 = {1{`RANDOM}};
  lengths_230 = _RAND_807[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_808 = {1{`RANDOM}};
  lengths_231 = _RAND_808[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_809 = {1{`RANDOM}};
  lengths_232 = _RAND_809[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_810 = {1{`RANDOM}};
  lengths_233 = _RAND_810[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_811 = {1{`RANDOM}};
  lengths_234 = _RAND_811[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_812 = {1{`RANDOM}};
  lengths_235 = _RAND_812[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_813 = {1{`RANDOM}};
  lengths_236 = _RAND_813[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_814 = {1{`RANDOM}};
  lengths_237 = _RAND_814[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_815 = {1{`RANDOM}};
  lengths_238 = _RAND_815[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_816 = {1{`RANDOM}};
  lengths_239 = _RAND_816[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_817 = {1{`RANDOM}};
  lengths_240 = _RAND_817[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_818 = {1{`RANDOM}};
  lengths_241 = _RAND_818[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_819 = {1{`RANDOM}};
  lengths_242 = _RAND_819[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_820 = {1{`RANDOM}};
  lengths_243 = _RAND_820[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_821 = {1{`RANDOM}};
  lengths_244 = _RAND_821[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_822 = {1{`RANDOM}};
  lengths_245 = _RAND_822[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_823 = {1{`RANDOM}};
  lengths_246 = _RAND_823[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_824 = {1{`RANDOM}};
  lengths_247 = _RAND_824[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_825 = {1{`RANDOM}};
  lengths_248 = _RAND_825[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_826 = {1{`RANDOM}};
  lengths_249 = _RAND_826[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_827 = {1{`RANDOM}};
  lengths_250 = _RAND_827[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_828 = {1{`RANDOM}};
  lengths_251 = _RAND_828[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_829 = {1{`RANDOM}};
  lengths_252 = _RAND_829[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_830 = {1{`RANDOM}};
  lengths_253 = _RAND_830[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_831 = {1{`RANDOM}};
  lengths_254 = _RAND_831[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_832 = {1{`RANDOM}};
  lengths_255 = _RAND_832[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_833 = {1{`RANDOM}};
  lengthsOut_0 = _RAND_833[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_834 = {1{`RANDOM}};
  lengthsOut_1 = _RAND_834[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_835 = {1{`RANDOM}};
  lengthsOut_2 = _RAND_835[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_836 = {1{`RANDOM}};
  lengthsOut_3 = _RAND_836[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_837 = {1{`RANDOM}};
  lengthsOut_4 = _RAND_837[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_838 = {1{`RANDOM}};
  lengthsOut_5 = _RAND_838[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_839 = {1{`RANDOM}};
  lengthsOut_6 = _RAND_839[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_840 = {1{`RANDOM}};
  lengthsOut_7 = _RAND_840[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_841 = {1{`RANDOM}};
  lengthsOut_8 = _RAND_841[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_842 = {1{`RANDOM}};
  lengthsOut_9 = _RAND_842[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_843 = {1{`RANDOM}};
  lengthsOut_10 = _RAND_843[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_844 = {1{`RANDOM}};
  lengthsOut_11 = _RAND_844[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_845 = {1{`RANDOM}};
  lengthsOut_12 = _RAND_845[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_846 = {1{`RANDOM}};
  lengthsOut_13 = _RAND_846[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_847 = {1{`RANDOM}};
  lengthsOut_14 = _RAND_847[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_848 = {1{`RANDOM}};
  lengthsOut_15 = _RAND_848[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_849 = {1{`RANDOM}};
  lengthsOut_16 = _RAND_849[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_850 = {1{`RANDOM}};
  lengthsOut_17 = _RAND_850[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_851 = {1{`RANDOM}};
  lengthsOut_18 = _RAND_851[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_852 = {1{`RANDOM}};
  lengthsOut_19 = _RAND_852[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_853 = {1{`RANDOM}};
  lengthsOut_20 = _RAND_853[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_854 = {1{`RANDOM}};
  lengthsOut_21 = _RAND_854[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_855 = {1{`RANDOM}};
  lengthsOut_22 = _RAND_855[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_856 = {1{`RANDOM}};
  lengthsOut_23 = _RAND_856[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_857 = {1{`RANDOM}};
  lengthsOut_24 = _RAND_857[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_858 = {1{`RANDOM}};
  lengthsOut_25 = _RAND_858[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_859 = {1{`RANDOM}};
  lengthsOut_26 = _RAND_859[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_860 = {1{`RANDOM}};
  lengthsOut_27 = _RAND_860[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_861 = {1{`RANDOM}};
  lengthsOut_28 = _RAND_861[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_862 = {1{`RANDOM}};
  lengthsOut_29 = _RAND_862[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_863 = {1{`RANDOM}};
  lengthsOut_30 = _RAND_863[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_864 = {1{`RANDOM}};
  lengthsOut_31 = _RAND_864[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_865 = {1{`RANDOM}};
  lengthsOut_32 = _RAND_865[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_866 = {1{`RANDOM}};
  lengthsOut_33 = _RAND_866[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_867 = {1{`RANDOM}};
  lengthsOut_34 = _RAND_867[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_868 = {1{`RANDOM}};
  lengthsOut_35 = _RAND_868[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_869 = {1{`RANDOM}};
  lengthsOut_36 = _RAND_869[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_870 = {1{`RANDOM}};
  lengthsOut_37 = _RAND_870[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_871 = {1{`RANDOM}};
  lengthsOut_38 = _RAND_871[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_872 = {1{`RANDOM}};
  lengthsOut_39 = _RAND_872[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_873 = {1{`RANDOM}};
  lengthsOut_40 = _RAND_873[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_874 = {1{`RANDOM}};
  lengthsOut_41 = _RAND_874[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_875 = {1{`RANDOM}};
  lengthsOut_42 = _RAND_875[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_876 = {1{`RANDOM}};
  lengthsOut_43 = _RAND_876[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_877 = {1{`RANDOM}};
  lengthsOut_44 = _RAND_877[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_878 = {1{`RANDOM}};
  lengthsOut_45 = _RAND_878[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_879 = {1{`RANDOM}};
  lengthsOut_46 = _RAND_879[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_880 = {1{`RANDOM}};
  lengthsOut_47 = _RAND_880[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_881 = {1{`RANDOM}};
  lengthsOut_48 = _RAND_881[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_882 = {1{`RANDOM}};
  lengthsOut_49 = _RAND_882[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_883 = {1{`RANDOM}};
  lengthsOut_50 = _RAND_883[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_884 = {1{`RANDOM}};
  lengthsOut_51 = _RAND_884[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_885 = {1{`RANDOM}};
  lengthsOut_52 = _RAND_885[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_886 = {1{`RANDOM}};
  lengthsOut_53 = _RAND_886[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_887 = {1{`RANDOM}};
  lengthsOut_54 = _RAND_887[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_888 = {1{`RANDOM}};
  lengthsOut_55 = _RAND_888[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_889 = {1{`RANDOM}};
  lengthsOut_56 = _RAND_889[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_890 = {1{`RANDOM}};
  lengthsOut_57 = _RAND_890[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_891 = {1{`RANDOM}};
  lengthsOut_58 = _RAND_891[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_892 = {1{`RANDOM}};
  lengthsOut_59 = _RAND_892[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_893 = {1{`RANDOM}};
  lengthsOut_60 = _RAND_893[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_894 = {1{`RANDOM}};
  lengthsOut_61 = _RAND_894[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_895 = {1{`RANDOM}};
  lengthsOut_62 = _RAND_895[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_896 = {1{`RANDOM}};
  lengthsOut_63 = _RAND_896[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_897 = {1{`RANDOM}};
  lengthsOut_64 = _RAND_897[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_898 = {1{`RANDOM}};
  lengthsOut_65 = _RAND_898[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_899 = {1{`RANDOM}};
  lengthsOut_66 = _RAND_899[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_900 = {1{`RANDOM}};
  lengthsOut_67 = _RAND_900[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_901 = {1{`RANDOM}};
  lengthsOut_68 = _RAND_901[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_902 = {1{`RANDOM}};
  lengthsOut_69 = _RAND_902[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_903 = {1{`RANDOM}};
  lengthsOut_70 = _RAND_903[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_904 = {1{`RANDOM}};
  lengthsOut_71 = _RAND_904[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_905 = {1{`RANDOM}};
  lengthsOut_72 = _RAND_905[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_906 = {1{`RANDOM}};
  lengthsOut_73 = _RAND_906[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_907 = {1{`RANDOM}};
  lengthsOut_74 = _RAND_907[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_908 = {1{`RANDOM}};
  lengthsOut_75 = _RAND_908[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_909 = {1{`RANDOM}};
  lengthsOut_76 = _RAND_909[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_910 = {1{`RANDOM}};
  lengthsOut_77 = _RAND_910[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_911 = {1{`RANDOM}};
  lengthsOut_78 = _RAND_911[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_912 = {1{`RANDOM}};
  lengthsOut_79 = _RAND_912[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_913 = {1{`RANDOM}};
  lengthsOut_80 = _RAND_913[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_914 = {1{`RANDOM}};
  lengthsOut_81 = _RAND_914[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_915 = {1{`RANDOM}};
  lengthsOut_82 = _RAND_915[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_916 = {1{`RANDOM}};
  lengthsOut_83 = _RAND_916[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_917 = {1{`RANDOM}};
  lengthsOut_84 = _RAND_917[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_918 = {1{`RANDOM}};
  lengthsOut_85 = _RAND_918[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_919 = {1{`RANDOM}};
  lengthsOut_86 = _RAND_919[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_920 = {1{`RANDOM}};
  lengthsOut_87 = _RAND_920[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_921 = {1{`RANDOM}};
  lengthsOut_88 = _RAND_921[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_922 = {1{`RANDOM}};
  lengthsOut_89 = _RAND_922[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_923 = {1{`RANDOM}};
  lengthsOut_90 = _RAND_923[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_924 = {1{`RANDOM}};
  lengthsOut_91 = _RAND_924[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_925 = {1{`RANDOM}};
  lengthsOut_92 = _RAND_925[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_926 = {1{`RANDOM}};
  lengthsOut_93 = _RAND_926[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_927 = {1{`RANDOM}};
  lengthsOut_94 = _RAND_927[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_928 = {1{`RANDOM}};
  lengthsOut_95 = _RAND_928[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_929 = {1{`RANDOM}};
  lengthsOut_96 = _RAND_929[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_930 = {1{`RANDOM}};
  lengthsOut_97 = _RAND_930[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_931 = {1{`RANDOM}};
  lengthsOut_98 = _RAND_931[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_932 = {1{`RANDOM}};
  lengthsOut_99 = _RAND_932[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_933 = {1{`RANDOM}};
  lengthsOut_100 = _RAND_933[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_934 = {1{`RANDOM}};
  lengthsOut_101 = _RAND_934[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_935 = {1{`RANDOM}};
  lengthsOut_102 = _RAND_935[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_936 = {1{`RANDOM}};
  lengthsOut_103 = _RAND_936[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_937 = {1{`RANDOM}};
  lengthsOut_104 = _RAND_937[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_938 = {1{`RANDOM}};
  lengthsOut_105 = _RAND_938[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_939 = {1{`RANDOM}};
  lengthsOut_106 = _RAND_939[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_940 = {1{`RANDOM}};
  lengthsOut_107 = _RAND_940[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_941 = {1{`RANDOM}};
  lengthsOut_108 = _RAND_941[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_942 = {1{`RANDOM}};
  lengthsOut_109 = _RAND_942[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_943 = {1{`RANDOM}};
  lengthsOut_110 = _RAND_943[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_944 = {1{`RANDOM}};
  lengthsOut_111 = _RAND_944[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_945 = {1{`RANDOM}};
  lengthsOut_112 = _RAND_945[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_946 = {1{`RANDOM}};
  lengthsOut_113 = _RAND_946[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_947 = {1{`RANDOM}};
  lengthsOut_114 = _RAND_947[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_948 = {1{`RANDOM}};
  lengthsOut_115 = _RAND_948[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_949 = {1{`RANDOM}};
  lengthsOut_116 = _RAND_949[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_950 = {1{`RANDOM}};
  lengthsOut_117 = _RAND_950[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_951 = {1{`RANDOM}};
  lengthsOut_118 = _RAND_951[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_952 = {1{`RANDOM}};
  lengthsOut_119 = _RAND_952[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_953 = {1{`RANDOM}};
  lengthsOut_120 = _RAND_953[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_954 = {1{`RANDOM}};
  lengthsOut_121 = _RAND_954[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_955 = {1{`RANDOM}};
  lengthsOut_122 = _RAND_955[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_956 = {1{`RANDOM}};
  lengthsOut_123 = _RAND_956[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_957 = {1{`RANDOM}};
  lengthsOut_124 = _RAND_957[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_958 = {1{`RANDOM}};
  lengthsOut_125 = _RAND_958[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_959 = {1{`RANDOM}};
  lengthsOut_126 = _RAND_959[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_960 = {1{`RANDOM}};
  lengthsOut_127 = _RAND_960[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_961 = {1{`RANDOM}};
  lengthsOut_128 = _RAND_961[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_962 = {1{`RANDOM}};
  lengthsOut_129 = _RAND_962[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_963 = {1{`RANDOM}};
  lengthsOut_130 = _RAND_963[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_964 = {1{`RANDOM}};
  lengthsOut_131 = _RAND_964[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_965 = {1{`RANDOM}};
  lengthsOut_132 = _RAND_965[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_966 = {1{`RANDOM}};
  lengthsOut_133 = _RAND_966[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_967 = {1{`RANDOM}};
  lengthsOut_134 = _RAND_967[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_968 = {1{`RANDOM}};
  lengthsOut_135 = _RAND_968[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_969 = {1{`RANDOM}};
  lengthsOut_136 = _RAND_969[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_970 = {1{`RANDOM}};
  lengthsOut_137 = _RAND_970[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_971 = {1{`RANDOM}};
  lengthsOut_138 = _RAND_971[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_972 = {1{`RANDOM}};
  lengthsOut_139 = _RAND_972[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_973 = {1{`RANDOM}};
  lengthsOut_140 = _RAND_973[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_974 = {1{`RANDOM}};
  lengthsOut_141 = _RAND_974[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_975 = {1{`RANDOM}};
  lengthsOut_142 = _RAND_975[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_976 = {1{`RANDOM}};
  lengthsOut_143 = _RAND_976[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_977 = {1{`RANDOM}};
  lengthsOut_144 = _RAND_977[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_978 = {1{`RANDOM}};
  lengthsOut_145 = _RAND_978[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_979 = {1{`RANDOM}};
  lengthsOut_146 = _RAND_979[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_980 = {1{`RANDOM}};
  lengthsOut_147 = _RAND_980[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_981 = {1{`RANDOM}};
  lengthsOut_148 = _RAND_981[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_982 = {1{`RANDOM}};
  lengthsOut_149 = _RAND_982[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_983 = {1{`RANDOM}};
  lengthsOut_150 = _RAND_983[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_984 = {1{`RANDOM}};
  lengthsOut_151 = _RAND_984[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_985 = {1{`RANDOM}};
  lengthsOut_152 = _RAND_985[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_986 = {1{`RANDOM}};
  lengthsOut_153 = _RAND_986[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_987 = {1{`RANDOM}};
  lengthsOut_154 = _RAND_987[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_988 = {1{`RANDOM}};
  lengthsOut_155 = _RAND_988[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_989 = {1{`RANDOM}};
  lengthsOut_156 = _RAND_989[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_990 = {1{`RANDOM}};
  lengthsOut_157 = _RAND_990[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_991 = {1{`RANDOM}};
  lengthsOut_158 = _RAND_991[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_992 = {1{`RANDOM}};
  lengthsOut_159 = _RAND_992[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_993 = {1{`RANDOM}};
  lengthsOut_160 = _RAND_993[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_994 = {1{`RANDOM}};
  lengthsOut_161 = _RAND_994[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_995 = {1{`RANDOM}};
  lengthsOut_162 = _RAND_995[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_996 = {1{`RANDOM}};
  lengthsOut_163 = _RAND_996[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_997 = {1{`RANDOM}};
  lengthsOut_164 = _RAND_997[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_998 = {1{`RANDOM}};
  lengthsOut_165 = _RAND_998[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_999 = {1{`RANDOM}};
  lengthsOut_166 = _RAND_999[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1000 = {1{`RANDOM}};
  lengthsOut_167 = _RAND_1000[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1001 = {1{`RANDOM}};
  lengthsOut_168 = _RAND_1001[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1002 = {1{`RANDOM}};
  lengthsOut_169 = _RAND_1002[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1003 = {1{`RANDOM}};
  lengthsOut_170 = _RAND_1003[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1004 = {1{`RANDOM}};
  lengthsOut_171 = _RAND_1004[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1005 = {1{`RANDOM}};
  lengthsOut_172 = _RAND_1005[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1006 = {1{`RANDOM}};
  lengthsOut_173 = _RAND_1006[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1007 = {1{`RANDOM}};
  lengthsOut_174 = _RAND_1007[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1008 = {1{`RANDOM}};
  lengthsOut_175 = _RAND_1008[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1009 = {1{`RANDOM}};
  lengthsOut_176 = _RAND_1009[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1010 = {1{`RANDOM}};
  lengthsOut_177 = _RAND_1010[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1011 = {1{`RANDOM}};
  lengthsOut_178 = _RAND_1011[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1012 = {1{`RANDOM}};
  lengthsOut_179 = _RAND_1012[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1013 = {1{`RANDOM}};
  lengthsOut_180 = _RAND_1013[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1014 = {1{`RANDOM}};
  lengthsOut_181 = _RAND_1014[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1015 = {1{`RANDOM}};
  lengthsOut_182 = _RAND_1015[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1016 = {1{`RANDOM}};
  lengthsOut_183 = _RAND_1016[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1017 = {1{`RANDOM}};
  lengthsOut_184 = _RAND_1017[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1018 = {1{`RANDOM}};
  lengthsOut_185 = _RAND_1018[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1019 = {1{`RANDOM}};
  lengthsOut_186 = _RAND_1019[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1020 = {1{`RANDOM}};
  lengthsOut_187 = _RAND_1020[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1021 = {1{`RANDOM}};
  lengthsOut_188 = _RAND_1021[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1022 = {1{`RANDOM}};
  lengthsOut_189 = _RAND_1022[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1023 = {1{`RANDOM}};
  lengthsOut_190 = _RAND_1023[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1024 = {1{`RANDOM}};
  lengthsOut_191 = _RAND_1024[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1025 = {1{`RANDOM}};
  lengthsOut_192 = _RAND_1025[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1026 = {1{`RANDOM}};
  lengthsOut_193 = _RAND_1026[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1027 = {1{`RANDOM}};
  lengthsOut_194 = _RAND_1027[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1028 = {1{`RANDOM}};
  lengthsOut_195 = _RAND_1028[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1029 = {1{`RANDOM}};
  lengthsOut_196 = _RAND_1029[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1030 = {1{`RANDOM}};
  lengthsOut_197 = _RAND_1030[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1031 = {1{`RANDOM}};
  lengthsOut_198 = _RAND_1031[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1032 = {1{`RANDOM}};
  lengthsOut_199 = _RAND_1032[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1033 = {1{`RANDOM}};
  lengthsOut_200 = _RAND_1033[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1034 = {1{`RANDOM}};
  lengthsOut_201 = _RAND_1034[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1035 = {1{`RANDOM}};
  lengthsOut_202 = _RAND_1035[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1036 = {1{`RANDOM}};
  lengthsOut_203 = _RAND_1036[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1037 = {1{`RANDOM}};
  lengthsOut_204 = _RAND_1037[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1038 = {1{`RANDOM}};
  lengthsOut_205 = _RAND_1038[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1039 = {1{`RANDOM}};
  lengthsOut_206 = _RAND_1039[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1040 = {1{`RANDOM}};
  lengthsOut_207 = _RAND_1040[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1041 = {1{`RANDOM}};
  lengthsOut_208 = _RAND_1041[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1042 = {1{`RANDOM}};
  lengthsOut_209 = _RAND_1042[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1043 = {1{`RANDOM}};
  lengthsOut_210 = _RAND_1043[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1044 = {1{`RANDOM}};
  lengthsOut_211 = _RAND_1044[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1045 = {1{`RANDOM}};
  lengthsOut_212 = _RAND_1045[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1046 = {1{`RANDOM}};
  lengthsOut_213 = _RAND_1046[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1047 = {1{`RANDOM}};
  lengthsOut_214 = _RAND_1047[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1048 = {1{`RANDOM}};
  lengthsOut_215 = _RAND_1048[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1049 = {1{`RANDOM}};
  lengthsOut_216 = _RAND_1049[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1050 = {1{`RANDOM}};
  lengthsOut_217 = _RAND_1050[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1051 = {1{`RANDOM}};
  lengthsOut_218 = _RAND_1051[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1052 = {1{`RANDOM}};
  lengthsOut_219 = _RAND_1052[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1053 = {1{`RANDOM}};
  lengthsOut_220 = _RAND_1053[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1054 = {1{`RANDOM}};
  lengthsOut_221 = _RAND_1054[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1055 = {1{`RANDOM}};
  lengthsOut_222 = _RAND_1055[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1056 = {1{`RANDOM}};
  lengthsOut_223 = _RAND_1056[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1057 = {1{`RANDOM}};
  lengthsOut_224 = _RAND_1057[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1058 = {1{`RANDOM}};
  lengthsOut_225 = _RAND_1058[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1059 = {1{`RANDOM}};
  lengthsOut_226 = _RAND_1059[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1060 = {1{`RANDOM}};
  lengthsOut_227 = _RAND_1060[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1061 = {1{`RANDOM}};
  lengthsOut_228 = _RAND_1061[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1062 = {1{`RANDOM}};
  lengthsOut_229 = _RAND_1062[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1063 = {1{`RANDOM}};
  lengthsOut_230 = _RAND_1063[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1064 = {1{`RANDOM}};
  lengthsOut_231 = _RAND_1064[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1065 = {1{`RANDOM}};
  lengthsOut_232 = _RAND_1065[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1066 = {1{`RANDOM}};
  lengthsOut_233 = _RAND_1066[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1067 = {1{`RANDOM}};
  lengthsOut_234 = _RAND_1067[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1068 = {1{`RANDOM}};
  lengthsOut_235 = _RAND_1068[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1069 = {1{`RANDOM}};
  lengthsOut_236 = _RAND_1069[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1070 = {1{`RANDOM}};
  lengthsOut_237 = _RAND_1070[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1071 = {1{`RANDOM}};
  lengthsOut_238 = _RAND_1071[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1072 = {1{`RANDOM}};
  lengthsOut_239 = _RAND_1072[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1073 = {1{`RANDOM}};
  lengthsOut_240 = _RAND_1073[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1074 = {1{`RANDOM}};
  lengthsOut_241 = _RAND_1074[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1075 = {1{`RANDOM}};
  lengthsOut_242 = _RAND_1075[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1076 = {1{`RANDOM}};
  lengthsOut_243 = _RAND_1076[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1077 = {1{`RANDOM}};
  lengthsOut_244 = _RAND_1077[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1078 = {1{`RANDOM}};
  lengthsOut_245 = _RAND_1078[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1079 = {1{`RANDOM}};
  lengthsOut_246 = _RAND_1079[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1080 = {1{`RANDOM}};
  lengthsOut_247 = _RAND_1080[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1081 = {1{`RANDOM}};
  lengthsOut_248 = _RAND_1081[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1082 = {1{`RANDOM}};
  lengthsOut_249 = _RAND_1082[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1083 = {1{`RANDOM}};
  lengthsOut_250 = _RAND_1083[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1084 = {1{`RANDOM}};
  lengthsOut_251 = _RAND_1084[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1085 = {1{`RANDOM}};
  lengthsOut_252 = _RAND_1085[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1086 = {1{`RANDOM}};
  lengthsOut_253 = _RAND_1086[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1087 = {1{`RANDOM}};
  lengthsOut_254 = _RAND_1087[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1088 = {1{`RANDOM}};
  lengthsOut_255 = _RAND_1088[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1089 = {1{`RANDOM}};
  characterIndex = _RAND_1089[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1090 = {1{`RANDOM}};
  nodes = _RAND_1090[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1091 = {1{`RANDOM}};
  characterDepth = _RAND_1091[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1092 = {1{`RANDOM}};
  codeword = _RAND_1092[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1093 = {1{`RANDOM}};
  escapeCodeword = _RAND_1093[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1094 = {1{`RANDOM}};
  escapeCharacterLength = _RAND_1094[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T_6) begin
      if (io_start) begin
        state <= 2'h1;
      end
    end else if (_T_9) begin
      if (_T_29) begin
        state <= 2'h2;
      end
    end else if (_T_30) begin
      if (_T_29) begin
        state <= 2'h3;
      end
    end else if (_T_65) begin
      state <= 2'h0;
    end
    if (reset) begin
      charactersIn_0 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_0 <= io_inputs_charactersOut_0;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h0 == _T_12[4:0]) begin
            if (5'h1f == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_31;
            end else if (5'h1e == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_30;
            end else if (5'h1d == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_29;
            end else if (5'h1c == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_28;
            end else if (5'h1b == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_27;
            end else if (5'h1a == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_26;
            end else if (5'h19 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_25;
            end else if (5'h18 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_24;
            end else if (5'h17 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_23;
            end else if (5'h16 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_22;
            end else if (5'h15 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_21;
            end else if (5'h14 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_20;
            end else if (5'h13 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_19;
            end else if (5'h12 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_18;
            end else if (5'h11 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_17;
            end else if (5'h10 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_16;
            end else if (5'hf == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_15;
            end else if (5'he == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_14;
            end else if (5'hd == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_13;
            end else if (5'hc == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_12;
            end else if (5'hb == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_11;
            end else if (5'ha == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_10;
            end else if (5'h9 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_9;
            end else if (5'h8 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_8;
            end else if (5'h7 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_7;
            end else if (5'h6 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_6;
            end else if (5'h5 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_5;
            end else if (5'h4 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_4;
            end else if (5'h3 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_3;
            end else if (5'h2 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_2;
            end else if (5'h1 == characterIndex[4:0]) begin
              charactersIn_0 <= charactersIn_1;
            end
          end else if (5'h0 == characterIndex[4:0]) begin
            if (5'h1f == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_31;
            end else if (5'h1e == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_30;
            end else if (5'h1d == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_29;
            end else if (5'h1c == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_28;
            end else if (5'h1b == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_27;
            end else if (5'h1a == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_26;
            end else if (5'h19 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_25;
            end else if (5'h18 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_24;
            end else if (5'h17 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_23;
            end else if (5'h16 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_22;
            end else if (5'h15 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_21;
            end else if (5'h14 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_20;
            end else if (5'h13 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_19;
            end else if (5'h12 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_18;
            end else if (5'h11 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_17;
            end else if (5'h10 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_16;
            end else if (5'hf == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_15;
            end else if (5'he == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_14;
            end else if (5'hd == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_13;
            end else if (5'hc == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_12;
            end else if (5'hb == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_11;
            end else if (5'ha == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_10;
            end else if (5'h9 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_9;
            end else if (5'h8 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_8;
            end else if (5'h7 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_7;
            end else if (5'h6 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_6;
            end else if (5'h5 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_5;
            end else if (5'h4 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_4;
            end else if (5'h3 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_3;
            end else if (5'h2 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_2;
            end else if (5'h1 == _T_12[4:0]) begin
              charactersIn_0 <= charactersIn_1;
            end
          end
        end
      end
    end
    if (reset) begin
      charactersIn_1 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_1 <= io_inputs_charactersOut_1;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h1 == _T_12[4:0]) begin
            if (5'h1f == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_31;
            end else if (5'h1e == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_30;
            end else if (5'h1d == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_29;
            end else if (5'h1c == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_28;
            end else if (5'h1b == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_27;
            end else if (5'h1a == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_26;
            end else if (5'h19 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_25;
            end else if (5'h18 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_24;
            end else if (5'h17 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_23;
            end else if (5'h16 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_22;
            end else if (5'h15 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_21;
            end else if (5'h14 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_20;
            end else if (5'h13 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_19;
            end else if (5'h12 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_18;
            end else if (5'h11 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_17;
            end else if (5'h10 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_16;
            end else if (5'hf == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_15;
            end else if (5'he == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_14;
            end else if (5'hd == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_13;
            end else if (5'hc == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_12;
            end else if (5'hb == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_11;
            end else if (5'ha == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_10;
            end else if (5'h9 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_9;
            end else if (5'h8 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_8;
            end else if (5'h7 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_7;
            end else if (5'h6 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_6;
            end else if (5'h5 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_5;
            end else if (5'h4 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_4;
            end else if (5'h3 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_3;
            end else if (5'h2 == characterIndex[4:0]) begin
              charactersIn_1 <= charactersIn_2;
            end else if (!(5'h1 == characterIndex[4:0])) begin
              charactersIn_1 <= charactersIn_0;
            end
          end else if (5'h1 == characterIndex[4:0]) begin
            if (5'h1f == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_31;
            end else if (5'h1e == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_30;
            end else if (5'h1d == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_29;
            end else if (5'h1c == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_28;
            end else if (5'h1b == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_27;
            end else if (5'h1a == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_26;
            end else if (5'h19 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_25;
            end else if (5'h18 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_24;
            end else if (5'h17 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_23;
            end else if (5'h16 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_22;
            end else if (5'h15 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_21;
            end else if (5'h14 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_20;
            end else if (5'h13 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_19;
            end else if (5'h12 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_18;
            end else if (5'h11 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_17;
            end else if (5'h10 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_16;
            end else if (5'hf == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_15;
            end else if (5'he == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_14;
            end else if (5'hd == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_13;
            end else if (5'hc == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_12;
            end else if (5'hb == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_11;
            end else if (5'ha == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_10;
            end else if (5'h9 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_9;
            end else if (5'h8 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_8;
            end else if (5'h7 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_7;
            end else if (5'h6 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_6;
            end else if (5'h5 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_5;
            end else if (5'h4 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_4;
            end else if (5'h3 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_3;
            end else if (5'h2 == _T_12[4:0]) begin
              charactersIn_1 <= charactersIn_2;
            end else if (!(5'h1 == _T_12[4:0])) begin
              charactersIn_1 <= charactersIn_0;
            end
          end
        end
      end
    end
    if (reset) begin
      charactersIn_2 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_2 <= io_inputs_charactersOut_2;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h2 == _T_12[4:0]) begin
            if (5'h1f == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_31;
            end else if (5'h1e == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_30;
            end else if (5'h1d == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_29;
            end else if (5'h1c == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_28;
            end else if (5'h1b == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_27;
            end else if (5'h1a == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_26;
            end else if (5'h19 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_25;
            end else if (5'h18 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_24;
            end else if (5'h17 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_23;
            end else if (5'h16 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_22;
            end else if (5'h15 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_21;
            end else if (5'h14 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_20;
            end else if (5'h13 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_19;
            end else if (5'h12 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_18;
            end else if (5'h11 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_17;
            end else if (5'h10 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_16;
            end else if (5'hf == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_15;
            end else if (5'he == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_14;
            end else if (5'hd == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_13;
            end else if (5'hc == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_12;
            end else if (5'hb == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_11;
            end else if (5'ha == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_10;
            end else if (5'h9 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_9;
            end else if (5'h8 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_8;
            end else if (5'h7 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_7;
            end else if (5'h6 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_6;
            end else if (5'h5 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_5;
            end else if (5'h4 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_4;
            end else if (5'h3 == characterIndex[4:0]) begin
              charactersIn_2 <= charactersIn_3;
            end else if (!(5'h2 == characterIndex[4:0])) begin
              if (5'h1 == characterIndex[4:0]) begin
                charactersIn_2 <= charactersIn_1;
              end else begin
                charactersIn_2 <= charactersIn_0;
              end
            end
          end else if (5'h2 == characterIndex[4:0]) begin
            if (5'h1f == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_31;
            end else if (5'h1e == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_30;
            end else if (5'h1d == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_29;
            end else if (5'h1c == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_28;
            end else if (5'h1b == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_27;
            end else if (5'h1a == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_26;
            end else if (5'h19 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_25;
            end else if (5'h18 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_24;
            end else if (5'h17 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_23;
            end else if (5'h16 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_22;
            end else if (5'h15 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_21;
            end else if (5'h14 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_20;
            end else if (5'h13 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_19;
            end else if (5'h12 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_18;
            end else if (5'h11 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_17;
            end else if (5'h10 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_16;
            end else if (5'hf == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_15;
            end else if (5'he == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_14;
            end else if (5'hd == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_13;
            end else if (5'hc == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_12;
            end else if (5'hb == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_11;
            end else if (5'ha == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_10;
            end else if (5'h9 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_9;
            end else if (5'h8 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_8;
            end else if (5'h7 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_7;
            end else if (5'h6 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_6;
            end else if (5'h5 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_5;
            end else if (5'h4 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_4;
            end else if (5'h3 == _T_12[4:0]) begin
              charactersIn_2 <= charactersIn_3;
            end else if (!(5'h2 == _T_12[4:0])) begin
              if (5'h1 == _T_12[4:0]) begin
                charactersIn_2 <= charactersIn_1;
              end else begin
                charactersIn_2 <= charactersIn_0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      charactersIn_3 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_3 <= io_inputs_charactersOut_3;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h3 == _T_12[4:0]) begin
            if (5'h1f == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_31;
            end else if (5'h1e == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_30;
            end else if (5'h1d == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_29;
            end else if (5'h1c == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_28;
            end else if (5'h1b == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_27;
            end else if (5'h1a == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_26;
            end else if (5'h19 == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_25;
            end else if (5'h18 == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_24;
            end else if (5'h17 == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_23;
            end else if (5'h16 == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_22;
            end else if (5'h15 == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_21;
            end else if (5'h14 == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_20;
            end else if (5'h13 == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_19;
            end else if (5'h12 == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_18;
            end else if (5'h11 == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_17;
            end else if (5'h10 == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_16;
            end else if (5'hf == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_15;
            end else if (5'he == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_14;
            end else if (5'hd == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_13;
            end else if (5'hc == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_12;
            end else if (5'hb == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_11;
            end else if (5'ha == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_10;
            end else if (5'h9 == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_9;
            end else if (5'h8 == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_8;
            end else if (5'h7 == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_7;
            end else if (5'h6 == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_6;
            end else if (5'h5 == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_5;
            end else if (5'h4 == characterIndex[4:0]) begin
              charactersIn_3 <= charactersIn_4;
            end else if (!(5'h3 == characterIndex[4:0])) begin
              if (5'h2 == characterIndex[4:0]) begin
                charactersIn_3 <= charactersIn_2;
              end else if (5'h1 == characterIndex[4:0]) begin
                charactersIn_3 <= charactersIn_1;
              end else begin
                charactersIn_3 <= charactersIn_0;
              end
            end
          end else if (5'h3 == characterIndex[4:0]) begin
            if (5'h1f == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_31;
            end else if (5'h1e == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_30;
            end else if (5'h1d == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_29;
            end else if (5'h1c == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_28;
            end else if (5'h1b == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_27;
            end else if (5'h1a == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_26;
            end else if (5'h19 == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_25;
            end else if (5'h18 == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_24;
            end else if (5'h17 == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_23;
            end else if (5'h16 == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_22;
            end else if (5'h15 == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_21;
            end else if (5'h14 == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_20;
            end else if (5'h13 == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_19;
            end else if (5'h12 == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_18;
            end else if (5'h11 == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_17;
            end else if (5'h10 == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_16;
            end else if (5'hf == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_15;
            end else if (5'he == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_14;
            end else if (5'hd == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_13;
            end else if (5'hc == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_12;
            end else if (5'hb == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_11;
            end else if (5'ha == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_10;
            end else if (5'h9 == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_9;
            end else if (5'h8 == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_8;
            end else if (5'h7 == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_7;
            end else if (5'h6 == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_6;
            end else if (5'h5 == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_5;
            end else if (5'h4 == _T_12[4:0]) begin
              charactersIn_3 <= charactersIn_4;
            end else if (!(5'h3 == _T_12[4:0])) begin
              if (5'h2 == _T_12[4:0]) begin
                charactersIn_3 <= charactersIn_2;
              end else if (5'h1 == _T_12[4:0]) begin
                charactersIn_3 <= charactersIn_1;
              end else begin
                charactersIn_3 <= charactersIn_0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      charactersIn_4 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_4 <= io_inputs_charactersOut_4;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h4 == _T_12[4:0]) begin
            charactersIn_4 <= _GEN_182;
          end else if (5'h4 == characterIndex[4:0]) begin
            charactersIn_4 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_5 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_5 <= io_inputs_charactersOut_5;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h5 == _T_12[4:0]) begin
            charactersIn_5 <= _GEN_182;
          end else if (5'h5 == characterIndex[4:0]) begin
            charactersIn_5 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_6 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_6 <= io_inputs_charactersOut_6;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h6 == _T_12[4:0]) begin
            charactersIn_6 <= _GEN_182;
          end else if (5'h6 == characterIndex[4:0]) begin
            charactersIn_6 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_7 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_7 <= io_inputs_charactersOut_7;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h7 == _T_12[4:0]) begin
            charactersIn_7 <= _GEN_182;
          end else if (5'h7 == characterIndex[4:0]) begin
            charactersIn_7 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_8 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_8 <= io_inputs_charactersOut_8;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h8 == _T_12[4:0]) begin
            charactersIn_8 <= _GEN_182;
          end else if (5'h8 == characterIndex[4:0]) begin
            charactersIn_8 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_9 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_9 <= io_inputs_charactersOut_9;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h9 == _T_12[4:0]) begin
            charactersIn_9 <= _GEN_182;
          end else if (5'h9 == characterIndex[4:0]) begin
            charactersIn_9 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_10 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_10 <= io_inputs_charactersOut_10;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'ha == _T_12[4:0]) begin
            charactersIn_10 <= _GEN_182;
          end else if (5'ha == characterIndex[4:0]) begin
            charactersIn_10 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_11 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_11 <= io_inputs_charactersOut_11;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'hb == _T_12[4:0]) begin
            charactersIn_11 <= _GEN_182;
          end else if (5'hb == characterIndex[4:0]) begin
            charactersIn_11 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_12 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_12 <= io_inputs_charactersOut_12;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'hc == _T_12[4:0]) begin
            charactersIn_12 <= _GEN_182;
          end else if (5'hc == characterIndex[4:0]) begin
            charactersIn_12 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_13 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_13 <= io_inputs_charactersOut_13;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'hd == _T_12[4:0]) begin
            charactersIn_13 <= _GEN_182;
          end else if (5'hd == characterIndex[4:0]) begin
            charactersIn_13 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_14 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_14 <= io_inputs_charactersOut_14;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'he == _T_12[4:0]) begin
            charactersIn_14 <= _GEN_182;
          end else if (5'he == characterIndex[4:0]) begin
            charactersIn_14 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_15 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_15 <= io_inputs_charactersOut_15;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'hf == _T_12[4:0]) begin
            charactersIn_15 <= _GEN_182;
          end else if (5'hf == characterIndex[4:0]) begin
            charactersIn_15 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_16 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_16 <= io_inputs_charactersOut_16;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h10 == _T_12[4:0]) begin
            charactersIn_16 <= _GEN_182;
          end else if (5'h10 == characterIndex[4:0]) begin
            charactersIn_16 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_17 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_17 <= io_inputs_charactersOut_17;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h11 == _T_12[4:0]) begin
            charactersIn_17 <= _GEN_182;
          end else if (5'h11 == characterIndex[4:0]) begin
            charactersIn_17 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_18 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_18 <= io_inputs_charactersOut_18;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h12 == _T_12[4:0]) begin
            charactersIn_18 <= _GEN_182;
          end else if (5'h12 == characterIndex[4:0]) begin
            charactersIn_18 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_19 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_19 <= io_inputs_charactersOut_19;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h13 == _T_12[4:0]) begin
            charactersIn_19 <= _GEN_182;
          end else if (5'h13 == characterIndex[4:0]) begin
            charactersIn_19 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_20 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_20 <= io_inputs_charactersOut_20;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h14 == _T_12[4:0]) begin
            charactersIn_20 <= _GEN_182;
          end else if (5'h14 == characterIndex[4:0]) begin
            charactersIn_20 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_21 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_21 <= io_inputs_charactersOut_21;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h15 == _T_12[4:0]) begin
            charactersIn_21 <= _GEN_182;
          end else if (5'h15 == characterIndex[4:0]) begin
            charactersIn_21 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_22 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_22 <= io_inputs_charactersOut_22;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h16 == _T_12[4:0]) begin
            charactersIn_22 <= _GEN_182;
          end else if (5'h16 == characterIndex[4:0]) begin
            charactersIn_22 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_23 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_23 <= io_inputs_charactersOut_23;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h17 == _T_12[4:0]) begin
            charactersIn_23 <= _GEN_182;
          end else if (5'h17 == characterIndex[4:0]) begin
            charactersIn_23 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_24 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_24 <= io_inputs_charactersOut_24;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h18 == _T_12[4:0]) begin
            charactersIn_24 <= _GEN_182;
          end else if (5'h18 == characterIndex[4:0]) begin
            charactersIn_24 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_25 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_25 <= io_inputs_charactersOut_25;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h19 == _T_12[4:0]) begin
            charactersIn_25 <= _GEN_182;
          end else if (5'h19 == characterIndex[4:0]) begin
            charactersIn_25 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_26 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_26 <= io_inputs_charactersOut_26;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h1a == _T_12[4:0]) begin
            charactersIn_26 <= _GEN_182;
          end else if (5'h1a == characterIndex[4:0]) begin
            charactersIn_26 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_27 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_27 <= io_inputs_charactersOut_27;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h1b == _T_12[4:0]) begin
            charactersIn_27 <= _GEN_182;
          end else if (5'h1b == characterIndex[4:0]) begin
            charactersIn_27 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_28 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_28 <= io_inputs_charactersOut_28;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h1c == _T_12[4:0]) begin
            charactersIn_28 <= _GEN_182;
          end else if (5'h1c == characterIndex[4:0]) begin
            charactersIn_28 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_29 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_29 <= io_inputs_charactersOut_29;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h1d == _T_12[4:0]) begin
            charactersIn_29 <= _GEN_182;
          end else if (5'h1d == characterIndex[4:0]) begin
            charactersIn_29 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_30 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_30 <= io_inputs_charactersOut_30;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h1e == _T_12[4:0]) begin
            charactersIn_30 <= _GEN_182;
          end else if (5'h1e == characterIndex[4:0]) begin
            charactersIn_30 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      charactersIn_31 <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        charactersIn_31 <= io_inputs_charactersOut_31;
      end
    end else if (_T_9) begin
      if (_T_14) begin
        if (_T_16) begin
          if (5'h1f == _T_12[4:0]) begin
            charactersIn_31 <= _GEN_182;
          end else if (5'h1f == characterIndex[4:0]) begin
            charactersIn_31 <= _GEN_246;
          end
        end
      end
    end
    if (reset) begin
      depths_0 <= 4'h0;
    end else begin
      depths_0 <= _GEN_7784[3:0];
    end
    if (reset) begin
      depths_1 <= 4'h0;
    end else begin
      depths_1 <= _GEN_7785[3:0];
    end
    if (reset) begin
      depths_2 <= 4'h0;
    end else begin
      depths_2 <= _GEN_7786[3:0];
    end
    if (reset) begin
      depths_3 <= 4'h0;
    end else begin
      depths_3 <= _GEN_7787[3:0];
    end
    if (reset) begin
      depths_4 <= 4'h0;
    end else begin
      depths_4 <= _GEN_7788[3:0];
    end
    if (reset) begin
      depths_5 <= 4'h0;
    end else begin
      depths_5 <= _GEN_7789[3:0];
    end
    if (reset) begin
      depths_6 <= 4'h0;
    end else begin
      depths_6 <= _GEN_7790[3:0];
    end
    if (reset) begin
      depths_7 <= 4'h0;
    end else begin
      depths_7 <= _GEN_7791[3:0];
    end
    if (reset) begin
      depths_8 <= 4'h0;
    end else begin
      depths_8 <= _GEN_7792[3:0];
    end
    if (reset) begin
      depths_9 <= 4'h0;
    end else begin
      depths_9 <= _GEN_7793[3:0];
    end
    if (reset) begin
      depths_10 <= 4'h0;
    end else begin
      depths_10 <= _GEN_7794[3:0];
    end
    if (reset) begin
      depths_11 <= 4'h0;
    end else begin
      depths_11 <= _GEN_7795[3:0];
    end
    if (reset) begin
      depths_12 <= 4'h0;
    end else begin
      depths_12 <= _GEN_7796[3:0];
    end
    if (reset) begin
      depths_13 <= 4'h0;
    end else begin
      depths_13 <= _GEN_7797[3:0];
    end
    if (reset) begin
      depths_14 <= 4'h0;
    end else begin
      depths_14 <= _GEN_7798[3:0];
    end
    if (reset) begin
      depths_15 <= 4'h0;
    end else begin
      depths_15 <= _GEN_7799[3:0];
    end
    if (reset) begin
      depths_16 <= 4'h0;
    end else begin
      depths_16 <= _GEN_7800[3:0];
    end
    if (reset) begin
      depths_17 <= 4'h0;
    end else begin
      depths_17 <= _GEN_7801[3:0];
    end
    if (reset) begin
      depths_18 <= 4'h0;
    end else begin
      depths_18 <= _GEN_7802[3:0];
    end
    if (reset) begin
      depths_19 <= 4'h0;
    end else begin
      depths_19 <= _GEN_7803[3:0];
    end
    if (reset) begin
      depths_20 <= 4'h0;
    end else begin
      depths_20 <= _GEN_7804[3:0];
    end
    if (reset) begin
      depths_21 <= 4'h0;
    end else begin
      depths_21 <= _GEN_7805[3:0];
    end
    if (reset) begin
      depths_22 <= 4'h0;
    end else begin
      depths_22 <= _GEN_7806[3:0];
    end
    if (reset) begin
      depths_23 <= 4'h0;
    end else begin
      depths_23 <= _GEN_7807[3:0];
    end
    if (reset) begin
      depths_24 <= 4'h0;
    end else begin
      depths_24 <= _GEN_7808[3:0];
    end
    if (reset) begin
      depths_25 <= 4'h0;
    end else begin
      depths_25 <= _GEN_7809[3:0];
    end
    if (reset) begin
      depths_26 <= 4'h0;
    end else begin
      depths_26 <= _GEN_7810[3:0];
    end
    if (reset) begin
      depths_27 <= 4'h0;
    end else begin
      depths_27 <= _GEN_7811[3:0];
    end
    if (reset) begin
      depths_28 <= 4'h0;
    end else begin
      depths_28 <= _GEN_7812[3:0];
    end
    if (reset) begin
      depths_29 <= 4'h0;
    end else begin
      depths_29 <= _GEN_7813[3:0];
    end
    if (reset) begin
      depths_30 <= 4'h0;
    end else begin
      depths_30 <= _GEN_7814[3:0];
    end
    if (reset) begin
      depths_31 <= 4'h0;
    end else begin
      depths_31 <= _GEN_7815[3:0];
    end
    if (reset) begin
      codewords_0 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h0 == _GEN_182[7:0]) begin
                codewords_0 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_1 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h1 == _GEN_182[7:0]) begin
                codewords_1 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_2 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h2 == _GEN_182[7:0]) begin
                codewords_2 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_3 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h3 == _GEN_182[7:0]) begin
                codewords_3 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_4 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h4 == _GEN_182[7:0]) begin
                codewords_4 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_5 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h5 == _GEN_182[7:0]) begin
                codewords_5 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_6 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h6 == _GEN_182[7:0]) begin
                codewords_6 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_7 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h7 == _GEN_182[7:0]) begin
                codewords_7 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_8 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h8 == _GEN_182[7:0]) begin
                codewords_8 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_9 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h9 == _GEN_182[7:0]) begin
                codewords_9 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_10 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha == _GEN_182[7:0]) begin
                codewords_10 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_11 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb == _GEN_182[7:0]) begin
                codewords_11 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_12 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc == _GEN_182[7:0]) begin
                codewords_12 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_13 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd == _GEN_182[7:0]) begin
                codewords_13 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_14 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he == _GEN_182[7:0]) begin
                codewords_14 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_15 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf == _GEN_182[7:0]) begin
                codewords_15 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_16 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h10 == _GEN_182[7:0]) begin
                codewords_16 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_17 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h11 == _GEN_182[7:0]) begin
                codewords_17 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_18 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h12 == _GEN_182[7:0]) begin
                codewords_18 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_19 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h13 == _GEN_182[7:0]) begin
                codewords_19 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_20 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h14 == _GEN_182[7:0]) begin
                codewords_20 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_21 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h15 == _GEN_182[7:0]) begin
                codewords_21 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_22 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h16 == _GEN_182[7:0]) begin
                codewords_22 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_23 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h17 == _GEN_182[7:0]) begin
                codewords_23 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_24 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h18 == _GEN_182[7:0]) begin
                codewords_24 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_25 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h19 == _GEN_182[7:0]) begin
                codewords_25 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_26 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h1a == _GEN_182[7:0]) begin
                codewords_26 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_27 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h1b == _GEN_182[7:0]) begin
                codewords_27 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_28 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h1c == _GEN_182[7:0]) begin
                codewords_28 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_29 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h1d == _GEN_182[7:0]) begin
                codewords_29 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_30 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h1e == _GEN_182[7:0]) begin
                codewords_30 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_31 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h1f == _GEN_182[7:0]) begin
                codewords_31 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_32 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h20 == _GEN_182[7:0]) begin
                codewords_32 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_33 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h21 == _GEN_182[7:0]) begin
                codewords_33 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_34 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h22 == _GEN_182[7:0]) begin
                codewords_34 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_35 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h23 == _GEN_182[7:0]) begin
                codewords_35 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_36 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h24 == _GEN_182[7:0]) begin
                codewords_36 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_37 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h25 == _GEN_182[7:0]) begin
                codewords_37 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_38 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h26 == _GEN_182[7:0]) begin
                codewords_38 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_39 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h27 == _GEN_182[7:0]) begin
                codewords_39 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_40 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h28 == _GEN_182[7:0]) begin
                codewords_40 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_41 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h29 == _GEN_182[7:0]) begin
                codewords_41 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_42 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h2a == _GEN_182[7:0]) begin
                codewords_42 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_43 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h2b == _GEN_182[7:0]) begin
                codewords_43 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_44 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h2c == _GEN_182[7:0]) begin
                codewords_44 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_45 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h2d == _GEN_182[7:0]) begin
                codewords_45 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_46 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h2e == _GEN_182[7:0]) begin
                codewords_46 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_47 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h2f == _GEN_182[7:0]) begin
                codewords_47 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_48 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h30 == _GEN_182[7:0]) begin
                codewords_48 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_49 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h31 == _GEN_182[7:0]) begin
                codewords_49 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_50 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h32 == _GEN_182[7:0]) begin
                codewords_50 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_51 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h33 == _GEN_182[7:0]) begin
                codewords_51 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_52 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h34 == _GEN_182[7:0]) begin
                codewords_52 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_53 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h35 == _GEN_182[7:0]) begin
                codewords_53 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_54 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h36 == _GEN_182[7:0]) begin
                codewords_54 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_55 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h37 == _GEN_182[7:0]) begin
                codewords_55 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_56 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h38 == _GEN_182[7:0]) begin
                codewords_56 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_57 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h39 == _GEN_182[7:0]) begin
                codewords_57 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_58 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h3a == _GEN_182[7:0]) begin
                codewords_58 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_59 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h3b == _GEN_182[7:0]) begin
                codewords_59 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_60 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h3c == _GEN_182[7:0]) begin
                codewords_60 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_61 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h3d == _GEN_182[7:0]) begin
                codewords_61 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_62 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h3e == _GEN_182[7:0]) begin
                codewords_62 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_63 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h3f == _GEN_182[7:0]) begin
                codewords_63 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_64 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h40 == _GEN_182[7:0]) begin
                codewords_64 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_65 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h41 == _GEN_182[7:0]) begin
                codewords_65 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_66 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h42 == _GEN_182[7:0]) begin
                codewords_66 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_67 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h43 == _GEN_182[7:0]) begin
                codewords_67 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_68 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h44 == _GEN_182[7:0]) begin
                codewords_68 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_69 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h45 == _GEN_182[7:0]) begin
                codewords_69 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_70 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h46 == _GEN_182[7:0]) begin
                codewords_70 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_71 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h47 == _GEN_182[7:0]) begin
                codewords_71 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_72 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h48 == _GEN_182[7:0]) begin
                codewords_72 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_73 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h49 == _GEN_182[7:0]) begin
                codewords_73 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_74 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h4a == _GEN_182[7:0]) begin
                codewords_74 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_75 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h4b == _GEN_182[7:0]) begin
                codewords_75 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_76 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h4c == _GEN_182[7:0]) begin
                codewords_76 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_77 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h4d == _GEN_182[7:0]) begin
                codewords_77 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_78 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h4e == _GEN_182[7:0]) begin
                codewords_78 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_79 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h4f == _GEN_182[7:0]) begin
                codewords_79 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_80 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h50 == _GEN_182[7:0]) begin
                codewords_80 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_81 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h51 == _GEN_182[7:0]) begin
                codewords_81 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_82 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h52 == _GEN_182[7:0]) begin
                codewords_82 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_83 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h53 == _GEN_182[7:0]) begin
                codewords_83 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_84 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h54 == _GEN_182[7:0]) begin
                codewords_84 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_85 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h55 == _GEN_182[7:0]) begin
                codewords_85 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_86 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h56 == _GEN_182[7:0]) begin
                codewords_86 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_87 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h57 == _GEN_182[7:0]) begin
                codewords_87 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_88 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h58 == _GEN_182[7:0]) begin
                codewords_88 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_89 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h59 == _GEN_182[7:0]) begin
                codewords_89 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_90 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h5a == _GEN_182[7:0]) begin
                codewords_90 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_91 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h5b == _GEN_182[7:0]) begin
                codewords_91 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_92 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h5c == _GEN_182[7:0]) begin
                codewords_92 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_93 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h5d == _GEN_182[7:0]) begin
                codewords_93 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_94 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h5e == _GEN_182[7:0]) begin
                codewords_94 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_95 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h5f == _GEN_182[7:0]) begin
                codewords_95 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_96 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h60 == _GEN_182[7:0]) begin
                codewords_96 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_97 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h61 == _GEN_182[7:0]) begin
                codewords_97 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_98 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h62 == _GEN_182[7:0]) begin
                codewords_98 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_99 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h63 == _GEN_182[7:0]) begin
                codewords_99 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_100 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h64 == _GEN_182[7:0]) begin
                codewords_100 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_101 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h65 == _GEN_182[7:0]) begin
                codewords_101 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_102 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h66 == _GEN_182[7:0]) begin
                codewords_102 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_103 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h67 == _GEN_182[7:0]) begin
                codewords_103 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_104 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h68 == _GEN_182[7:0]) begin
                codewords_104 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_105 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h69 == _GEN_182[7:0]) begin
                codewords_105 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_106 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h6a == _GEN_182[7:0]) begin
                codewords_106 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_107 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h6b == _GEN_182[7:0]) begin
                codewords_107 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_108 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h6c == _GEN_182[7:0]) begin
                codewords_108 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_109 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h6d == _GEN_182[7:0]) begin
                codewords_109 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_110 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h6e == _GEN_182[7:0]) begin
                codewords_110 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_111 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h6f == _GEN_182[7:0]) begin
                codewords_111 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_112 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h70 == _GEN_182[7:0]) begin
                codewords_112 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_113 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h71 == _GEN_182[7:0]) begin
                codewords_113 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_114 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h72 == _GEN_182[7:0]) begin
                codewords_114 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_115 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h73 == _GEN_182[7:0]) begin
                codewords_115 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_116 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h74 == _GEN_182[7:0]) begin
                codewords_116 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_117 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h75 == _GEN_182[7:0]) begin
                codewords_117 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_118 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h76 == _GEN_182[7:0]) begin
                codewords_118 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_119 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h77 == _GEN_182[7:0]) begin
                codewords_119 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_120 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h78 == _GEN_182[7:0]) begin
                codewords_120 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_121 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h79 == _GEN_182[7:0]) begin
                codewords_121 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_122 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h7a == _GEN_182[7:0]) begin
                codewords_122 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_123 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h7b == _GEN_182[7:0]) begin
                codewords_123 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_124 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h7c == _GEN_182[7:0]) begin
                codewords_124 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_125 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h7d == _GEN_182[7:0]) begin
                codewords_125 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_126 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h7e == _GEN_182[7:0]) begin
                codewords_126 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_127 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h7f == _GEN_182[7:0]) begin
                codewords_127 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_128 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h80 == _GEN_182[7:0]) begin
                codewords_128 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_129 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h81 == _GEN_182[7:0]) begin
                codewords_129 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_130 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h82 == _GEN_182[7:0]) begin
                codewords_130 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_131 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h83 == _GEN_182[7:0]) begin
                codewords_131 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_132 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h84 == _GEN_182[7:0]) begin
                codewords_132 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_133 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h85 == _GEN_182[7:0]) begin
                codewords_133 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_134 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h86 == _GEN_182[7:0]) begin
                codewords_134 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_135 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h87 == _GEN_182[7:0]) begin
                codewords_135 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_136 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h88 == _GEN_182[7:0]) begin
                codewords_136 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_137 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h89 == _GEN_182[7:0]) begin
                codewords_137 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_138 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h8a == _GEN_182[7:0]) begin
                codewords_138 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_139 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h8b == _GEN_182[7:0]) begin
                codewords_139 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_140 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h8c == _GEN_182[7:0]) begin
                codewords_140 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_141 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h8d == _GEN_182[7:0]) begin
                codewords_141 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_142 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h8e == _GEN_182[7:0]) begin
                codewords_142 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_143 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h8f == _GEN_182[7:0]) begin
                codewords_143 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_144 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h90 == _GEN_182[7:0]) begin
                codewords_144 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_145 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h91 == _GEN_182[7:0]) begin
                codewords_145 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_146 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h92 == _GEN_182[7:0]) begin
                codewords_146 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_147 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h93 == _GEN_182[7:0]) begin
                codewords_147 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_148 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h94 == _GEN_182[7:0]) begin
                codewords_148 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_149 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h95 == _GEN_182[7:0]) begin
                codewords_149 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_150 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h96 == _GEN_182[7:0]) begin
                codewords_150 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_151 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h97 == _GEN_182[7:0]) begin
                codewords_151 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_152 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h98 == _GEN_182[7:0]) begin
                codewords_152 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_153 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h99 == _GEN_182[7:0]) begin
                codewords_153 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_154 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h9a == _GEN_182[7:0]) begin
                codewords_154 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_155 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h9b == _GEN_182[7:0]) begin
                codewords_155 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_156 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h9c == _GEN_182[7:0]) begin
                codewords_156 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_157 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h9d == _GEN_182[7:0]) begin
                codewords_157 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_158 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h9e == _GEN_182[7:0]) begin
                codewords_158 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_159 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h9f == _GEN_182[7:0]) begin
                codewords_159 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_160 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha0 == _GEN_182[7:0]) begin
                codewords_160 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_161 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha1 == _GEN_182[7:0]) begin
                codewords_161 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_162 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha2 == _GEN_182[7:0]) begin
                codewords_162 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_163 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha3 == _GEN_182[7:0]) begin
                codewords_163 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_164 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha4 == _GEN_182[7:0]) begin
                codewords_164 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_165 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha5 == _GEN_182[7:0]) begin
                codewords_165 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_166 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha6 == _GEN_182[7:0]) begin
                codewords_166 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_167 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha7 == _GEN_182[7:0]) begin
                codewords_167 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_168 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha8 == _GEN_182[7:0]) begin
                codewords_168 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_169 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha9 == _GEN_182[7:0]) begin
                codewords_169 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_170 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'haa == _GEN_182[7:0]) begin
                codewords_170 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_171 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hab == _GEN_182[7:0]) begin
                codewords_171 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_172 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hac == _GEN_182[7:0]) begin
                codewords_172 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_173 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'had == _GEN_182[7:0]) begin
                codewords_173 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_174 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hae == _GEN_182[7:0]) begin
                codewords_174 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_175 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'haf == _GEN_182[7:0]) begin
                codewords_175 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_176 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb0 == _GEN_182[7:0]) begin
                codewords_176 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_177 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb1 == _GEN_182[7:0]) begin
                codewords_177 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_178 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb2 == _GEN_182[7:0]) begin
                codewords_178 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_179 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb3 == _GEN_182[7:0]) begin
                codewords_179 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_180 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb4 == _GEN_182[7:0]) begin
                codewords_180 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_181 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb5 == _GEN_182[7:0]) begin
                codewords_181 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_182 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb6 == _GEN_182[7:0]) begin
                codewords_182 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_183 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb7 == _GEN_182[7:0]) begin
                codewords_183 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_184 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb8 == _GEN_182[7:0]) begin
                codewords_184 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_185 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb9 == _GEN_182[7:0]) begin
                codewords_185 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_186 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hba == _GEN_182[7:0]) begin
                codewords_186 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_187 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hbb == _GEN_182[7:0]) begin
                codewords_187 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_188 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hbc == _GEN_182[7:0]) begin
                codewords_188 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_189 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hbd == _GEN_182[7:0]) begin
                codewords_189 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_190 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hbe == _GEN_182[7:0]) begin
                codewords_190 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_191 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hbf == _GEN_182[7:0]) begin
                codewords_191 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_192 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc0 == _GEN_182[7:0]) begin
                codewords_192 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_193 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc1 == _GEN_182[7:0]) begin
                codewords_193 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_194 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc2 == _GEN_182[7:0]) begin
                codewords_194 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_195 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc3 == _GEN_182[7:0]) begin
                codewords_195 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_196 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc4 == _GEN_182[7:0]) begin
                codewords_196 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_197 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc5 == _GEN_182[7:0]) begin
                codewords_197 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_198 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc6 == _GEN_182[7:0]) begin
                codewords_198 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_199 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc7 == _GEN_182[7:0]) begin
                codewords_199 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_200 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc8 == _GEN_182[7:0]) begin
                codewords_200 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_201 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc9 == _GEN_182[7:0]) begin
                codewords_201 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_202 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hca == _GEN_182[7:0]) begin
                codewords_202 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_203 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hcb == _GEN_182[7:0]) begin
                codewords_203 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_204 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hcc == _GEN_182[7:0]) begin
                codewords_204 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_205 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hcd == _GEN_182[7:0]) begin
                codewords_205 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_206 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hce == _GEN_182[7:0]) begin
                codewords_206 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_207 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hcf == _GEN_182[7:0]) begin
                codewords_207 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_208 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd0 == _GEN_182[7:0]) begin
                codewords_208 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_209 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd1 == _GEN_182[7:0]) begin
                codewords_209 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_210 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd2 == _GEN_182[7:0]) begin
                codewords_210 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_211 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd3 == _GEN_182[7:0]) begin
                codewords_211 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_212 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd4 == _GEN_182[7:0]) begin
                codewords_212 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_213 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd5 == _GEN_182[7:0]) begin
                codewords_213 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_214 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd6 == _GEN_182[7:0]) begin
                codewords_214 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_215 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd7 == _GEN_182[7:0]) begin
                codewords_215 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_216 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd8 == _GEN_182[7:0]) begin
                codewords_216 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_217 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd9 == _GEN_182[7:0]) begin
                codewords_217 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_218 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hda == _GEN_182[7:0]) begin
                codewords_218 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_219 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hdb == _GEN_182[7:0]) begin
                codewords_219 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_220 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hdc == _GEN_182[7:0]) begin
                codewords_220 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_221 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hdd == _GEN_182[7:0]) begin
                codewords_221 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_222 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hde == _GEN_182[7:0]) begin
                codewords_222 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_223 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hdf == _GEN_182[7:0]) begin
                codewords_223 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_224 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he0 == _GEN_182[7:0]) begin
                codewords_224 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_225 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he1 == _GEN_182[7:0]) begin
                codewords_225 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_226 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he2 == _GEN_182[7:0]) begin
                codewords_226 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_227 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he3 == _GEN_182[7:0]) begin
                codewords_227 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_228 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he4 == _GEN_182[7:0]) begin
                codewords_228 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_229 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he5 == _GEN_182[7:0]) begin
                codewords_229 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_230 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he6 == _GEN_182[7:0]) begin
                codewords_230 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_231 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he7 == _GEN_182[7:0]) begin
                codewords_231 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_232 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he8 == _GEN_182[7:0]) begin
                codewords_232 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_233 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he9 == _GEN_182[7:0]) begin
                codewords_233 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_234 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hea == _GEN_182[7:0]) begin
                codewords_234 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_235 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'heb == _GEN_182[7:0]) begin
                codewords_235 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_236 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hec == _GEN_182[7:0]) begin
                codewords_236 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_237 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hed == _GEN_182[7:0]) begin
                codewords_237 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_238 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hee == _GEN_182[7:0]) begin
                codewords_238 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_239 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hef == _GEN_182[7:0]) begin
                codewords_239 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_240 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf0 == _GEN_182[7:0]) begin
                codewords_240 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_241 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf1 == _GEN_182[7:0]) begin
                codewords_241 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_242 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf2 == _GEN_182[7:0]) begin
                codewords_242 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_243 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf3 == _GEN_182[7:0]) begin
                codewords_243 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_244 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf4 == _GEN_182[7:0]) begin
                codewords_244 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_245 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf5 == _GEN_182[7:0]) begin
                codewords_245 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_246 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf6 == _GEN_182[7:0]) begin
                codewords_246 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_247 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf7 == _GEN_182[7:0]) begin
                codewords_247 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_248 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf8 == _GEN_182[7:0]) begin
                codewords_248 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_249 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf9 == _GEN_182[7:0]) begin
                codewords_249 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_250 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hfa == _GEN_182[7:0]) begin
                codewords_250 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_251 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hfb == _GEN_182[7:0]) begin
                codewords_251 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_252 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hfc == _GEN_182[7:0]) begin
                codewords_252 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_253 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hfd == _GEN_182[7:0]) begin
                codewords_253 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_254 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hfe == _GEN_182[7:0]) begin
                codewords_254 <= codeword;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      codewords_255 <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hff == _GEN_182[7:0]) begin
                codewords_255 <= codeword;
              end
            end
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h0 == characterIndex) begin
              codewordsOut_0 <= _T_67;
            end
          end else if (8'h0 == characterIndex) begin
            codewordsOut_0 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h1 == characterIndex) begin
              codewordsOut_1 <= _T_67;
            end
          end else if (8'h1 == characterIndex) begin
            codewordsOut_1 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h2 == characterIndex) begin
              codewordsOut_2 <= _T_67;
            end
          end else if (8'h2 == characterIndex) begin
            codewordsOut_2 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h3 == characterIndex) begin
              codewordsOut_3 <= _T_67;
            end
          end else if (8'h3 == characterIndex) begin
            codewordsOut_3 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h4 == characterIndex) begin
              codewordsOut_4 <= _T_67;
            end
          end else if (8'h4 == characterIndex) begin
            codewordsOut_4 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h5 == characterIndex) begin
              codewordsOut_5 <= _T_67;
            end
          end else if (8'h5 == characterIndex) begin
            codewordsOut_5 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h6 == characterIndex) begin
              codewordsOut_6 <= _T_67;
            end
          end else if (8'h6 == characterIndex) begin
            codewordsOut_6 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h7 == characterIndex) begin
              codewordsOut_7 <= _T_67;
            end
          end else if (8'h7 == characterIndex) begin
            codewordsOut_7 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h8 == characterIndex) begin
              codewordsOut_8 <= _T_67;
            end
          end else if (8'h8 == characterIndex) begin
            codewordsOut_8 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h9 == characterIndex) begin
              codewordsOut_9 <= _T_67;
            end
          end else if (8'h9 == characterIndex) begin
            codewordsOut_9 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha == characterIndex) begin
              codewordsOut_10 <= _T_67;
            end
          end else if (8'ha == characterIndex) begin
            codewordsOut_10 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb == characterIndex) begin
              codewordsOut_11 <= _T_67;
            end
          end else if (8'hb == characterIndex) begin
            codewordsOut_11 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc == characterIndex) begin
              codewordsOut_12 <= _T_67;
            end
          end else if (8'hc == characterIndex) begin
            codewordsOut_12 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd == characterIndex) begin
              codewordsOut_13 <= _T_67;
            end
          end else if (8'hd == characterIndex) begin
            codewordsOut_13 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he == characterIndex) begin
              codewordsOut_14 <= _T_67;
            end
          end else if (8'he == characterIndex) begin
            codewordsOut_14 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf == characterIndex) begin
              codewordsOut_15 <= _T_67;
            end
          end else if (8'hf == characterIndex) begin
            codewordsOut_15 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h10 == characterIndex) begin
              codewordsOut_16 <= _T_67;
            end
          end else if (8'h10 == characterIndex) begin
            codewordsOut_16 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h11 == characterIndex) begin
              codewordsOut_17 <= _T_67;
            end
          end else if (8'h11 == characterIndex) begin
            codewordsOut_17 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h12 == characterIndex) begin
              codewordsOut_18 <= _T_67;
            end
          end else if (8'h12 == characterIndex) begin
            codewordsOut_18 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h13 == characterIndex) begin
              codewordsOut_19 <= _T_67;
            end
          end else if (8'h13 == characterIndex) begin
            codewordsOut_19 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h14 == characterIndex) begin
              codewordsOut_20 <= _T_67;
            end
          end else if (8'h14 == characterIndex) begin
            codewordsOut_20 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h15 == characterIndex) begin
              codewordsOut_21 <= _T_67;
            end
          end else if (8'h15 == characterIndex) begin
            codewordsOut_21 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h16 == characterIndex) begin
              codewordsOut_22 <= _T_67;
            end
          end else if (8'h16 == characterIndex) begin
            codewordsOut_22 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h17 == characterIndex) begin
              codewordsOut_23 <= _T_67;
            end
          end else if (8'h17 == characterIndex) begin
            codewordsOut_23 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h18 == characterIndex) begin
              codewordsOut_24 <= _T_67;
            end
          end else if (8'h18 == characterIndex) begin
            codewordsOut_24 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h19 == characterIndex) begin
              codewordsOut_25 <= _T_67;
            end
          end else if (8'h19 == characterIndex) begin
            codewordsOut_25 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h1a == characterIndex) begin
              codewordsOut_26 <= _T_67;
            end
          end else if (8'h1a == characterIndex) begin
            codewordsOut_26 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h1b == characterIndex) begin
              codewordsOut_27 <= _T_67;
            end
          end else if (8'h1b == characterIndex) begin
            codewordsOut_27 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h1c == characterIndex) begin
              codewordsOut_28 <= _T_67;
            end
          end else if (8'h1c == characterIndex) begin
            codewordsOut_28 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h1d == characterIndex) begin
              codewordsOut_29 <= _T_67;
            end
          end else if (8'h1d == characterIndex) begin
            codewordsOut_29 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h1e == characterIndex) begin
              codewordsOut_30 <= _T_67;
            end
          end else if (8'h1e == characterIndex) begin
            codewordsOut_30 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h1f == characterIndex) begin
              codewordsOut_31 <= _T_67;
            end
          end else if (8'h1f == characterIndex) begin
            codewordsOut_31 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h20 == characterIndex) begin
              codewordsOut_32 <= _T_67;
            end
          end else if (8'h20 == characterIndex) begin
            codewordsOut_32 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h21 == characterIndex) begin
              codewordsOut_33 <= _T_67;
            end
          end else if (8'h21 == characterIndex) begin
            codewordsOut_33 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h22 == characterIndex) begin
              codewordsOut_34 <= _T_67;
            end
          end else if (8'h22 == characterIndex) begin
            codewordsOut_34 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h23 == characterIndex) begin
              codewordsOut_35 <= _T_67;
            end
          end else if (8'h23 == characterIndex) begin
            codewordsOut_35 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h24 == characterIndex) begin
              codewordsOut_36 <= _T_67;
            end
          end else if (8'h24 == characterIndex) begin
            codewordsOut_36 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h25 == characterIndex) begin
              codewordsOut_37 <= _T_67;
            end
          end else if (8'h25 == characterIndex) begin
            codewordsOut_37 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h26 == characterIndex) begin
              codewordsOut_38 <= _T_67;
            end
          end else if (8'h26 == characterIndex) begin
            codewordsOut_38 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h27 == characterIndex) begin
              codewordsOut_39 <= _T_67;
            end
          end else if (8'h27 == characterIndex) begin
            codewordsOut_39 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h28 == characterIndex) begin
              codewordsOut_40 <= _T_67;
            end
          end else if (8'h28 == characterIndex) begin
            codewordsOut_40 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h29 == characterIndex) begin
              codewordsOut_41 <= _T_67;
            end
          end else if (8'h29 == characterIndex) begin
            codewordsOut_41 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h2a == characterIndex) begin
              codewordsOut_42 <= _T_67;
            end
          end else if (8'h2a == characterIndex) begin
            codewordsOut_42 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h2b == characterIndex) begin
              codewordsOut_43 <= _T_67;
            end
          end else if (8'h2b == characterIndex) begin
            codewordsOut_43 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h2c == characterIndex) begin
              codewordsOut_44 <= _T_67;
            end
          end else if (8'h2c == characterIndex) begin
            codewordsOut_44 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h2d == characterIndex) begin
              codewordsOut_45 <= _T_67;
            end
          end else if (8'h2d == characterIndex) begin
            codewordsOut_45 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h2e == characterIndex) begin
              codewordsOut_46 <= _T_67;
            end
          end else if (8'h2e == characterIndex) begin
            codewordsOut_46 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h2f == characterIndex) begin
              codewordsOut_47 <= _T_67;
            end
          end else if (8'h2f == characterIndex) begin
            codewordsOut_47 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h30 == characterIndex) begin
              codewordsOut_48 <= _T_67;
            end
          end else if (8'h30 == characterIndex) begin
            codewordsOut_48 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h31 == characterIndex) begin
              codewordsOut_49 <= _T_67;
            end
          end else if (8'h31 == characterIndex) begin
            codewordsOut_49 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h32 == characterIndex) begin
              codewordsOut_50 <= _T_67;
            end
          end else if (8'h32 == characterIndex) begin
            codewordsOut_50 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h33 == characterIndex) begin
              codewordsOut_51 <= _T_67;
            end
          end else if (8'h33 == characterIndex) begin
            codewordsOut_51 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h34 == characterIndex) begin
              codewordsOut_52 <= _T_67;
            end
          end else if (8'h34 == characterIndex) begin
            codewordsOut_52 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h35 == characterIndex) begin
              codewordsOut_53 <= _T_67;
            end
          end else if (8'h35 == characterIndex) begin
            codewordsOut_53 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h36 == characterIndex) begin
              codewordsOut_54 <= _T_67;
            end
          end else if (8'h36 == characterIndex) begin
            codewordsOut_54 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h37 == characterIndex) begin
              codewordsOut_55 <= _T_67;
            end
          end else if (8'h37 == characterIndex) begin
            codewordsOut_55 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h38 == characterIndex) begin
              codewordsOut_56 <= _T_67;
            end
          end else if (8'h38 == characterIndex) begin
            codewordsOut_56 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h39 == characterIndex) begin
              codewordsOut_57 <= _T_67;
            end
          end else if (8'h39 == characterIndex) begin
            codewordsOut_57 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h3a == characterIndex) begin
              codewordsOut_58 <= _T_67;
            end
          end else if (8'h3a == characterIndex) begin
            codewordsOut_58 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h3b == characterIndex) begin
              codewordsOut_59 <= _T_67;
            end
          end else if (8'h3b == characterIndex) begin
            codewordsOut_59 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h3c == characterIndex) begin
              codewordsOut_60 <= _T_67;
            end
          end else if (8'h3c == characterIndex) begin
            codewordsOut_60 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h3d == characterIndex) begin
              codewordsOut_61 <= _T_67;
            end
          end else if (8'h3d == characterIndex) begin
            codewordsOut_61 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h3e == characterIndex) begin
              codewordsOut_62 <= _T_67;
            end
          end else if (8'h3e == characterIndex) begin
            codewordsOut_62 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h3f == characterIndex) begin
              codewordsOut_63 <= _T_67;
            end
          end else if (8'h3f == characterIndex) begin
            codewordsOut_63 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h40 == characterIndex) begin
              codewordsOut_64 <= _T_67;
            end
          end else if (8'h40 == characterIndex) begin
            codewordsOut_64 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h41 == characterIndex) begin
              codewordsOut_65 <= _T_67;
            end
          end else if (8'h41 == characterIndex) begin
            codewordsOut_65 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h42 == characterIndex) begin
              codewordsOut_66 <= _T_67;
            end
          end else if (8'h42 == characterIndex) begin
            codewordsOut_66 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h43 == characterIndex) begin
              codewordsOut_67 <= _T_67;
            end
          end else if (8'h43 == characterIndex) begin
            codewordsOut_67 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h44 == characterIndex) begin
              codewordsOut_68 <= _T_67;
            end
          end else if (8'h44 == characterIndex) begin
            codewordsOut_68 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h45 == characterIndex) begin
              codewordsOut_69 <= _T_67;
            end
          end else if (8'h45 == characterIndex) begin
            codewordsOut_69 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h46 == characterIndex) begin
              codewordsOut_70 <= _T_67;
            end
          end else if (8'h46 == characterIndex) begin
            codewordsOut_70 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h47 == characterIndex) begin
              codewordsOut_71 <= _T_67;
            end
          end else if (8'h47 == characterIndex) begin
            codewordsOut_71 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h48 == characterIndex) begin
              codewordsOut_72 <= _T_67;
            end
          end else if (8'h48 == characterIndex) begin
            codewordsOut_72 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h49 == characterIndex) begin
              codewordsOut_73 <= _T_67;
            end
          end else if (8'h49 == characterIndex) begin
            codewordsOut_73 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h4a == characterIndex) begin
              codewordsOut_74 <= _T_67;
            end
          end else if (8'h4a == characterIndex) begin
            codewordsOut_74 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h4b == characterIndex) begin
              codewordsOut_75 <= _T_67;
            end
          end else if (8'h4b == characterIndex) begin
            codewordsOut_75 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h4c == characterIndex) begin
              codewordsOut_76 <= _T_67;
            end
          end else if (8'h4c == characterIndex) begin
            codewordsOut_76 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h4d == characterIndex) begin
              codewordsOut_77 <= _T_67;
            end
          end else if (8'h4d == characterIndex) begin
            codewordsOut_77 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h4e == characterIndex) begin
              codewordsOut_78 <= _T_67;
            end
          end else if (8'h4e == characterIndex) begin
            codewordsOut_78 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h4f == characterIndex) begin
              codewordsOut_79 <= _T_67;
            end
          end else if (8'h4f == characterIndex) begin
            codewordsOut_79 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h50 == characterIndex) begin
              codewordsOut_80 <= _T_67;
            end
          end else if (8'h50 == characterIndex) begin
            codewordsOut_80 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h51 == characterIndex) begin
              codewordsOut_81 <= _T_67;
            end
          end else if (8'h51 == characterIndex) begin
            codewordsOut_81 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h52 == characterIndex) begin
              codewordsOut_82 <= _T_67;
            end
          end else if (8'h52 == characterIndex) begin
            codewordsOut_82 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h53 == characterIndex) begin
              codewordsOut_83 <= _T_67;
            end
          end else if (8'h53 == characterIndex) begin
            codewordsOut_83 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h54 == characterIndex) begin
              codewordsOut_84 <= _T_67;
            end
          end else if (8'h54 == characterIndex) begin
            codewordsOut_84 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h55 == characterIndex) begin
              codewordsOut_85 <= _T_67;
            end
          end else if (8'h55 == characterIndex) begin
            codewordsOut_85 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h56 == characterIndex) begin
              codewordsOut_86 <= _T_67;
            end
          end else if (8'h56 == characterIndex) begin
            codewordsOut_86 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h57 == characterIndex) begin
              codewordsOut_87 <= _T_67;
            end
          end else if (8'h57 == characterIndex) begin
            codewordsOut_87 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h58 == characterIndex) begin
              codewordsOut_88 <= _T_67;
            end
          end else if (8'h58 == characterIndex) begin
            codewordsOut_88 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h59 == characterIndex) begin
              codewordsOut_89 <= _T_67;
            end
          end else if (8'h59 == characterIndex) begin
            codewordsOut_89 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h5a == characterIndex) begin
              codewordsOut_90 <= _T_67;
            end
          end else if (8'h5a == characterIndex) begin
            codewordsOut_90 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h5b == characterIndex) begin
              codewordsOut_91 <= _T_67;
            end
          end else if (8'h5b == characterIndex) begin
            codewordsOut_91 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h5c == characterIndex) begin
              codewordsOut_92 <= _T_67;
            end
          end else if (8'h5c == characterIndex) begin
            codewordsOut_92 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h5d == characterIndex) begin
              codewordsOut_93 <= _T_67;
            end
          end else if (8'h5d == characterIndex) begin
            codewordsOut_93 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h5e == characterIndex) begin
              codewordsOut_94 <= _T_67;
            end
          end else if (8'h5e == characterIndex) begin
            codewordsOut_94 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h5f == characterIndex) begin
              codewordsOut_95 <= _T_67;
            end
          end else if (8'h5f == characterIndex) begin
            codewordsOut_95 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h60 == characterIndex) begin
              codewordsOut_96 <= _T_67;
            end
          end else if (8'h60 == characterIndex) begin
            codewordsOut_96 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h61 == characterIndex) begin
              codewordsOut_97 <= _T_67;
            end
          end else if (8'h61 == characterIndex) begin
            codewordsOut_97 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h62 == characterIndex) begin
              codewordsOut_98 <= _T_67;
            end
          end else if (8'h62 == characterIndex) begin
            codewordsOut_98 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h63 == characterIndex) begin
              codewordsOut_99 <= _T_67;
            end
          end else if (8'h63 == characterIndex) begin
            codewordsOut_99 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h64 == characterIndex) begin
              codewordsOut_100 <= _T_67;
            end
          end else if (8'h64 == characterIndex) begin
            codewordsOut_100 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h65 == characterIndex) begin
              codewordsOut_101 <= _T_67;
            end
          end else if (8'h65 == characterIndex) begin
            codewordsOut_101 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h66 == characterIndex) begin
              codewordsOut_102 <= _T_67;
            end
          end else if (8'h66 == characterIndex) begin
            codewordsOut_102 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h67 == characterIndex) begin
              codewordsOut_103 <= _T_67;
            end
          end else if (8'h67 == characterIndex) begin
            codewordsOut_103 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h68 == characterIndex) begin
              codewordsOut_104 <= _T_67;
            end
          end else if (8'h68 == characterIndex) begin
            codewordsOut_104 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h69 == characterIndex) begin
              codewordsOut_105 <= _T_67;
            end
          end else if (8'h69 == characterIndex) begin
            codewordsOut_105 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h6a == characterIndex) begin
              codewordsOut_106 <= _T_67;
            end
          end else if (8'h6a == characterIndex) begin
            codewordsOut_106 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h6b == characterIndex) begin
              codewordsOut_107 <= _T_67;
            end
          end else if (8'h6b == characterIndex) begin
            codewordsOut_107 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h6c == characterIndex) begin
              codewordsOut_108 <= _T_67;
            end
          end else if (8'h6c == characterIndex) begin
            codewordsOut_108 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h6d == characterIndex) begin
              codewordsOut_109 <= _T_67;
            end
          end else if (8'h6d == characterIndex) begin
            codewordsOut_109 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h6e == characterIndex) begin
              codewordsOut_110 <= _T_67;
            end
          end else if (8'h6e == characterIndex) begin
            codewordsOut_110 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h6f == characterIndex) begin
              codewordsOut_111 <= _T_67;
            end
          end else if (8'h6f == characterIndex) begin
            codewordsOut_111 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h70 == characterIndex) begin
              codewordsOut_112 <= _T_67;
            end
          end else if (8'h70 == characterIndex) begin
            codewordsOut_112 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h71 == characterIndex) begin
              codewordsOut_113 <= _T_67;
            end
          end else if (8'h71 == characterIndex) begin
            codewordsOut_113 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h72 == characterIndex) begin
              codewordsOut_114 <= _T_67;
            end
          end else if (8'h72 == characterIndex) begin
            codewordsOut_114 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h73 == characterIndex) begin
              codewordsOut_115 <= _T_67;
            end
          end else if (8'h73 == characterIndex) begin
            codewordsOut_115 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h74 == characterIndex) begin
              codewordsOut_116 <= _T_67;
            end
          end else if (8'h74 == characterIndex) begin
            codewordsOut_116 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h75 == characterIndex) begin
              codewordsOut_117 <= _T_67;
            end
          end else if (8'h75 == characterIndex) begin
            codewordsOut_117 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h76 == characterIndex) begin
              codewordsOut_118 <= _T_67;
            end
          end else if (8'h76 == characterIndex) begin
            codewordsOut_118 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h77 == characterIndex) begin
              codewordsOut_119 <= _T_67;
            end
          end else if (8'h77 == characterIndex) begin
            codewordsOut_119 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h78 == characterIndex) begin
              codewordsOut_120 <= _T_67;
            end
          end else if (8'h78 == characterIndex) begin
            codewordsOut_120 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h79 == characterIndex) begin
              codewordsOut_121 <= _T_67;
            end
          end else if (8'h79 == characterIndex) begin
            codewordsOut_121 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h7a == characterIndex) begin
              codewordsOut_122 <= _T_67;
            end
          end else if (8'h7a == characterIndex) begin
            codewordsOut_122 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h7b == characterIndex) begin
              codewordsOut_123 <= _T_67;
            end
          end else if (8'h7b == characterIndex) begin
            codewordsOut_123 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h7c == characterIndex) begin
              codewordsOut_124 <= _T_67;
            end
          end else if (8'h7c == characterIndex) begin
            codewordsOut_124 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h7d == characterIndex) begin
              codewordsOut_125 <= _T_67;
            end
          end else if (8'h7d == characterIndex) begin
            codewordsOut_125 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h7e == characterIndex) begin
              codewordsOut_126 <= _T_67;
            end
          end else if (8'h7e == characterIndex) begin
            codewordsOut_126 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h7f == characterIndex) begin
              codewordsOut_127 <= _T_67;
            end
          end else if (8'h7f == characterIndex) begin
            codewordsOut_127 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h80 == characterIndex) begin
              codewordsOut_128 <= _T_67;
            end
          end else if (8'h80 == characterIndex) begin
            codewordsOut_128 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h81 == characterIndex) begin
              codewordsOut_129 <= _T_67;
            end
          end else if (8'h81 == characterIndex) begin
            codewordsOut_129 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h82 == characterIndex) begin
              codewordsOut_130 <= _T_67;
            end
          end else if (8'h82 == characterIndex) begin
            codewordsOut_130 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h83 == characterIndex) begin
              codewordsOut_131 <= _T_67;
            end
          end else if (8'h83 == characterIndex) begin
            codewordsOut_131 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h84 == characterIndex) begin
              codewordsOut_132 <= _T_67;
            end
          end else if (8'h84 == characterIndex) begin
            codewordsOut_132 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h85 == characterIndex) begin
              codewordsOut_133 <= _T_67;
            end
          end else if (8'h85 == characterIndex) begin
            codewordsOut_133 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h86 == characterIndex) begin
              codewordsOut_134 <= _T_67;
            end
          end else if (8'h86 == characterIndex) begin
            codewordsOut_134 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h87 == characterIndex) begin
              codewordsOut_135 <= _T_67;
            end
          end else if (8'h87 == characterIndex) begin
            codewordsOut_135 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h88 == characterIndex) begin
              codewordsOut_136 <= _T_67;
            end
          end else if (8'h88 == characterIndex) begin
            codewordsOut_136 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h89 == characterIndex) begin
              codewordsOut_137 <= _T_67;
            end
          end else if (8'h89 == characterIndex) begin
            codewordsOut_137 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h8a == characterIndex) begin
              codewordsOut_138 <= _T_67;
            end
          end else if (8'h8a == characterIndex) begin
            codewordsOut_138 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h8b == characterIndex) begin
              codewordsOut_139 <= _T_67;
            end
          end else if (8'h8b == characterIndex) begin
            codewordsOut_139 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h8c == characterIndex) begin
              codewordsOut_140 <= _T_67;
            end
          end else if (8'h8c == characterIndex) begin
            codewordsOut_140 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h8d == characterIndex) begin
              codewordsOut_141 <= _T_67;
            end
          end else if (8'h8d == characterIndex) begin
            codewordsOut_141 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h8e == characterIndex) begin
              codewordsOut_142 <= _T_67;
            end
          end else if (8'h8e == characterIndex) begin
            codewordsOut_142 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h8f == characterIndex) begin
              codewordsOut_143 <= _T_67;
            end
          end else if (8'h8f == characterIndex) begin
            codewordsOut_143 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h90 == characterIndex) begin
              codewordsOut_144 <= _T_67;
            end
          end else if (8'h90 == characterIndex) begin
            codewordsOut_144 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h91 == characterIndex) begin
              codewordsOut_145 <= _T_67;
            end
          end else if (8'h91 == characterIndex) begin
            codewordsOut_145 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h92 == characterIndex) begin
              codewordsOut_146 <= _T_67;
            end
          end else if (8'h92 == characterIndex) begin
            codewordsOut_146 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h93 == characterIndex) begin
              codewordsOut_147 <= _T_67;
            end
          end else if (8'h93 == characterIndex) begin
            codewordsOut_147 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h94 == characterIndex) begin
              codewordsOut_148 <= _T_67;
            end
          end else if (8'h94 == characterIndex) begin
            codewordsOut_148 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h95 == characterIndex) begin
              codewordsOut_149 <= _T_67;
            end
          end else if (8'h95 == characterIndex) begin
            codewordsOut_149 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h96 == characterIndex) begin
              codewordsOut_150 <= _T_67;
            end
          end else if (8'h96 == characterIndex) begin
            codewordsOut_150 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h97 == characterIndex) begin
              codewordsOut_151 <= _T_67;
            end
          end else if (8'h97 == characterIndex) begin
            codewordsOut_151 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h98 == characterIndex) begin
              codewordsOut_152 <= _T_67;
            end
          end else if (8'h98 == characterIndex) begin
            codewordsOut_152 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h99 == characterIndex) begin
              codewordsOut_153 <= _T_67;
            end
          end else if (8'h99 == characterIndex) begin
            codewordsOut_153 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h9a == characterIndex) begin
              codewordsOut_154 <= _T_67;
            end
          end else if (8'h9a == characterIndex) begin
            codewordsOut_154 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h9b == characterIndex) begin
              codewordsOut_155 <= _T_67;
            end
          end else if (8'h9b == characterIndex) begin
            codewordsOut_155 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h9c == characterIndex) begin
              codewordsOut_156 <= _T_67;
            end
          end else if (8'h9c == characterIndex) begin
            codewordsOut_156 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h9d == characterIndex) begin
              codewordsOut_157 <= _T_67;
            end
          end else if (8'h9d == characterIndex) begin
            codewordsOut_157 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h9e == characterIndex) begin
              codewordsOut_158 <= _T_67;
            end
          end else if (8'h9e == characterIndex) begin
            codewordsOut_158 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h9f == characterIndex) begin
              codewordsOut_159 <= _T_67;
            end
          end else if (8'h9f == characterIndex) begin
            codewordsOut_159 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha0 == characterIndex) begin
              codewordsOut_160 <= _T_67;
            end
          end else if (8'ha0 == characterIndex) begin
            codewordsOut_160 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha1 == characterIndex) begin
              codewordsOut_161 <= _T_67;
            end
          end else if (8'ha1 == characterIndex) begin
            codewordsOut_161 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha2 == characterIndex) begin
              codewordsOut_162 <= _T_67;
            end
          end else if (8'ha2 == characterIndex) begin
            codewordsOut_162 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha3 == characterIndex) begin
              codewordsOut_163 <= _T_67;
            end
          end else if (8'ha3 == characterIndex) begin
            codewordsOut_163 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha4 == characterIndex) begin
              codewordsOut_164 <= _T_67;
            end
          end else if (8'ha4 == characterIndex) begin
            codewordsOut_164 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha5 == characterIndex) begin
              codewordsOut_165 <= _T_67;
            end
          end else if (8'ha5 == characterIndex) begin
            codewordsOut_165 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha6 == characterIndex) begin
              codewordsOut_166 <= _T_67;
            end
          end else if (8'ha6 == characterIndex) begin
            codewordsOut_166 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha7 == characterIndex) begin
              codewordsOut_167 <= _T_67;
            end
          end else if (8'ha7 == characterIndex) begin
            codewordsOut_167 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha8 == characterIndex) begin
              codewordsOut_168 <= _T_67;
            end
          end else if (8'ha8 == characterIndex) begin
            codewordsOut_168 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha9 == characterIndex) begin
              codewordsOut_169 <= _T_67;
            end
          end else if (8'ha9 == characterIndex) begin
            codewordsOut_169 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'haa == characterIndex) begin
              codewordsOut_170 <= _T_67;
            end
          end else if (8'haa == characterIndex) begin
            codewordsOut_170 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hab == characterIndex) begin
              codewordsOut_171 <= _T_67;
            end
          end else if (8'hab == characterIndex) begin
            codewordsOut_171 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hac == characterIndex) begin
              codewordsOut_172 <= _T_67;
            end
          end else if (8'hac == characterIndex) begin
            codewordsOut_172 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'had == characterIndex) begin
              codewordsOut_173 <= _T_67;
            end
          end else if (8'had == characterIndex) begin
            codewordsOut_173 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hae == characterIndex) begin
              codewordsOut_174 <= _T_67;
            end
          end else if (8'hae == characterIndex) begin
            codewordsOut_174 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'haf == characterIndex) begin
              codewordsOut_175 <= _T_67;
            end
          end else if (8'haf == characterIndex) begin
            codewordsOut_175 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb0 == characterIndex) begin
              codewordsOut_176 <= _T_67;
            end
          end else if (8'hb0 == characterIndex) begin
            codewordsOut_176 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb1 == characterIndex) begin
              codewordsOut_177 <= _T_67;
            end
          end else if (8'hb1 == characterIndex) begin
            codewordsOut_177 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb2 == characterIndex) begin
              codewordsOut_178 <= _T_67;
            end
          end else if (8'hb2 == characterIndex) begin
            codewordsOut_178 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb3 == characterIndex) begin
              codewordsOut_179 <= _T_67;
            end
          end else if (8'hb3 == characterIndex) begin
            codewordsOut_179 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb4 == characterIndex) begin
              codewordsOut_180 <= _T_67;
            end
          end else if (8'hb4 == characterIndex) begin
            codewordsOut_180 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb5 == characterIndex) begin
              codewordsOut_181 <= _T_67;
            end
          end else if (8'hb5 == characterIndex) begin
            codewordsOut_181 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb6 == characterIndex) begin
              codewordsOut_182 <= _T_67;
            end
          end else if (8'hb6 == characterIndex) begin
            codewordsOut_182 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb7 == characterIndex) begin
              codewordsOut_183 <= _T_67;
            end
          end else if (8'hb7 == characterIndex) begin
            codewordsOut_183 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb8 == characterIndex) begin
              codewordsOut_184 <= _T_67;
            end
          end else if (8'hb8 == characterIndex) begin
            codewordsOut_184 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb9 == characterIndex) begin
              codewordsOut_185 <= _T_67;
            end
          end else if (8'hb9 == characterIndex) begin
            codewordsOut_185 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hba == characterIndex) begin
              codewordsOut_186 <= _T_67;
            end
          end else if (8'hba == characterIndex) begin
            codewordsOut_186 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hbb == characterIndex) begin
              codewordsOut_187 <= _T_67;
            end
          end else if (8'hbb == characterIndex) begin
            codewordsOut_187 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hbc == characterIndex) begin
              codewordsOut_188 <= _T_67;
            end
          end else if (8'hbc == characterIndex) begin
            codewordsOut_188 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hbd == characterIndex) begin
              codewordsOut_189 <= _T_67;
            end
          end else if (8'hbd == characterIndex) begin
            codewordsOut_189 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hbe == characterIndex) begin
              codewordsOut_190 <= _T_67;
            end
          end else if (8'hbe == characterIndex) begin
            codewordsOut_190 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hbf == characterIndex) begin
              codewordsOut_191 <= _T_67;
            end
          end else if (8'hbf == characterIndex) begin
            codewordsOut_191 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc0 == characterIndex) begin
              codewordsOut_192 <= _T_67;
            end
          end else if (8'hc0 == characterIndex) begin
            codewordsOut_192 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc1 == characterIndex) begin
              codewordsOut_193 <= _T_67;
            end
          end else if (8'hc1 == characterIndex) begin
            codewordsOut_193 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc2 == characterIndex) begin
              codewordsOut_194 <= _T_67;
            end
          end else if (8'hc2 == characterIndex) begin
            codewordsOut_194 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc3 == characterIndex) begin
              codewordsOut_195 <= _T_67;
            end
          end else if (8'hc3 == characterIndex) begin
            codewordsOut_195 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc4 == characterIndex) begin
              codewordsOut_196 <= _T_67;
            end
          end else if (8'hc4 == characterIndex) begin
            codewordsOut_196 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc5 == characterIndex) begin
              codewordsOut_197 <= _T_67;
            end
          end else if (8'hc5 == characterIndex) begin
            codewordsOut_197 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc6 == characterIndex) begin
              codewordsOut_198 <= _T_67;
            end
          end else if (8'hc6 == characterIndex) begin
            codewordsOut_198 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc7 == characterIndex) begin
              codewordsOut_199 <= _T_67;
            end
          end else if (8'hc7 == characterIndex) begin
            codewordsOut_199 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc8 == characterIndex) begin
              codewordsOut_200 <= _T_67;
            end
          end else if (8'hc8 == characterIndex) begin
            codewordsOut_200 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc9 == characterIndex) begin
              codewordsOut_201 <= _T_67;
            end
          end else if (8'hc9 == characterIndex) begin
            codewordsOut_201 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hca == characterIndex) begin
              codewordsOut_202 <= _T_67;
            end
          end else if (8'hca == characterIndex) begin
            codewordsOut_202 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hcb == characterIndex) begin
              codewordsOut_203 <= _T_67;
            end
          end else if (8'hcb == characterIndex) begin
            codewordsOut_203 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hcc == characterIndex) begin
              codewordsOut_204 <= _T_67;
            end
          end else if (8'hcc == characterIndex) begin
            codewordsOut_204 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hcd == characterIndex) begin
              codewordsOut_205 <= _T_67;
            end
          end else if (8'hcd == characterIndex) begin
            codewordsOut_205 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hce == characterIndex) begin
              codewordsOut_206 <= _T_67;
            end
          end else if (8'hce == characterIndex) begin
            codewordsOut_206 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hcf == characterIndex) begin
              codewordsOut_207 <= _T_67;
            end
          end else if (8'hcf == characterIndex) begin
            codewordsOut_207 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd0 == characterIndex) begin
              codewordsOut_208 <= _T_67;
            end
          end else if (8'hd0 == characterIndex) begin
            codewordsOut_208 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd1 == characterIndex) begin
              codewordsOut_209 <= _T_67;
            end
          end else if (8'hd1 == characterIndex) begin
            codewordsOut_209 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd2 == characterIndex) begin
              codewordsOut_210 <= _T_67;
            end
          end else if (8'hd2 == characterIndex) begin
            codewordsOut_210 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd3 == characterIndex) begin
              codewordsOut_211 <= _T_67;
            end
          end else if (8'hd3 == characterIndex) begin
            codewordsOut_211 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd4 == characterIndex) begin
              codewordsOut_212 <= _T_67;
            end
          end else if (8'hd4 == characterIndex) begin
            codewordsOut_212 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd5 == characterIndex) begin
              codewordsOut_213 <= _T_67;
            end
          end else if (8'hd5 == characterIndex) begin
            codewordsOut_213 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd6 == characterIndex) begin
              codewordsOut_214 <= _T_67;
            end
          end else if (8'hd6 == characterIndex) begin
            codewordsOut_214 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd7 == characterIndex) begin
              codewordsOut_215 <= _T_67;
            end
          end else if (8'hd7 == characterIndex) begin
            codewordsOut_215 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd8 == characterIndex) begin
              codewordsOut_216 <= _T_67;
            end
          end else if (8'hd8 == characterIndex) begin
            codewordsOut_216 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd9 == characterIndex) begin
              codewordsOut_217 <= _T_67;
            end
          end else if (8'hd9 == characterIndex) begin
            codewordsOut_217 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hda == characterIndex) begin
              codewordsOut_218 <= _T_67;
            end
          end else if (8'hda == characterIndex) begin
            codewordsOut_218 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hdb == characterIndex) begin
              codewordsOut_219 <= _T_67;
            end
          end else if (8'hdb == characterIndex) begin
            codewordsOut_219 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hdc == characterIndex) begin
              codewordsOut_220 <= _T_67;
            end
          end else if (8'hdc == characterIndex) begin
            codewordsOut_220 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hdd == characterIndex) begin
              codewordsOut_221 <= _T_67;
            end
          end else if (8'hdd == characterIndex) begin
            codewordsOut_221 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hde == characterIndex) begin
              codewordsOut_222 <= _T_67;
            end
          end else if (8'hde == characterIndex) begin
            codewordsOut_222 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hdf == characterIndex) begin
              codewordsOut_223 <= _T_67;
            end
          end else if (8'hdf == characterIndex) begin
            codewordsOut_223 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he0 == characterIndex) begin
              codewordsOut_224 <= _T_67;
            end
          end else if (8'he0 == characterIndex) begin
            codewordsOut_224 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he1 == characterIndex) begin
              codewordsOut_225 <= _T_67;
            end
          end else if (8'he1 == characterIndex) begin
            codewordsOut_225 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he2 == characterIndex) begin
              codewordsOut_226 <= _T_67;
            end
          end else if (8'he2 == characterIndex) begin
            codewordsOut_226 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he3 == characterIndex) begin
              codewordsOut_227 <= _T_67;
            end
          end else if (8'he3 == characterIndex) begin
            codewordsOut_227 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he4 == characterIndex) begin
              codewordsOut_228 <= _T_67;
            end
          end else if (8'he4 == characterIndex) begin
            codewordsOut_228 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he5 == characterIndex) begin
              codewordsOut_229 <= _T_67;
            end
          end else if (8'he5 == characterIndex) begin
            codewordsOut_229 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he6 == characterIndex) begin
              codewordsOut_230 <= _T_67;
            end
          end else if (8'he6 == characterIndex) begin
            codewordsOut_230 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he7 == characterIndex) begin
              codewordsOut_231 <= _T_67;
            end
          end else if (8'he7 == characterIndex) begin
            codewordsOut_231 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he8 == characterIndex) begin
              codewordsOut_232 <= _T_67;
            end
          end else if (8'he8 == characterIndex) begin
            codewordsOut_232 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he9 == characterIndex) begin
              codewordsOut_233 <= _T_67;
            end
          end else if (8'he9 == characterIndex) begin
            codewordsOut_233 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hea == characterIndex) begin
              codewordsOut_234 <= _T_67;
            end
          end else if (8'hea == characterIndex) begin
            codewordsOut_234 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'heb == characterIndex) begin
              codewordsOut_235 <= _T_67;
            end
          end else if (8'heb == characterIndex) begin
            codewordsOut_235 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hec == characterIndex) begin
              codewordsOut_236 <= _T_67;
            end
          end else if (8'hec == characterIndex) begin
            codewordsOut_236 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hed == characterIndex) begin
              codewordsOut_237 <= _T_67;
            end
          end else if (8'hed == characterIndex) begin
            codewordsOut_237 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hee == characterIndex) begin
              codewordsOut_238 <= _T_67;
            end
          end else if (8'hee == characterIndex) begin
            codewordsOut_238 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hef == characterIndex) begin
              codewordsOut_239 <= _T_67;
            end
          end else if (8'hef == characterIndex) begin
            codewordsOut_239 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf0 == characterIndex) begin
              codewordsOut_240 <= _T_67;
            end
          end else if (8'hf0 == characterIndex) begin
            codewordsOut_240 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf1 == characterIndex) begin
              codewordsOut_241 <= _T_67;
            end
          end else if (8'hf1 == characterIndex) begin
            codewordsOut_241 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf2 == characterIndex) begin
              codewordsOut_242 <= _T_67;
            end
          end else if (8'hf2 == characterIndex) begin
            codewordsOut_242 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf3 == characterIndex) begin
              codewordsOut_243 <= _T_67;
            end
          end else if (8'hf3 == characterIndex) begin
            codewordsOut_243 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf4 == characterIndex) begin
              codewordsOut_244 <= _T_67;
            end
          end else if (8'hf4 == characterIndex) begin
            codewordsOut_244 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf5 == characterIndex) begin
              codewordsOut_245 <= _T_67;
            end
          end else if (8'hf5 == characterIndex) begin
            codewordsOut_245 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf6 == characterIndex) begin
              codewordsOut_246 <= _T_67;
            end
          end else if (8'hf6 == characterIndex) begin
            codewordsOut_246 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf7 == characterIndex) begin
              codewordsOut_247 <= _T_67;
            end
          end else if (8'hf7 == characterIndex) begin
            codewordsOut_247 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf8 == characterIndex) begin
              codewordsOut_248 <= _T_67;
            end
          end else if (8'hf8 == characterIndex) begin
            codewordsOut_248 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf9 == characterIndex) begin
              codewordsOut_249 <= _T_67;
            end
          end else if (8'hf9 == characterIndex) begin
            codewordsOut_249 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hfa == characterIndex) begin
              codewordsOut_250 <= _T_67;
            end
          end else if (8'hfa == characterIndex) begin
            codewordsOut_250 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hfb == characterIndex) begin
              codewordsOut_251 <= _T_67;
            end
          end else if (8'hfb == characterIndex) begin
            codewordsOut_251 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hfc == characterIndex) begin
              codewordsOut_252 <= _T_67;
            end
          end else if (8'hfc == characterIndex) begin
            codewordsOut_252 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hfd == characterIndex) begin
              codewordsOut_253 <= _T_67;
            end
          end else if (8'hfd == characterIndex) begin
            codewordsOut_253 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hfe == characterIndex) begin
              codewordsOut_254 <= _T_67;
            end
          end else if (8'hfe == characterIndex) begin
            codewordsOut_254 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hff == characterIndex) begin
              codewordsOut_255 <= _T_67;
            end
          end else if (8'hff == characterIndex) begin
            codewordsOut_255 <= _codewordsOut_characterIndex_0;
          end
        end
      end
    end
    if (reset) begin
      lengths_0 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h0 == _GEN_182[7:0]) begin
                lengths_0 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_1 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h1 == _GEN_182[7:0]) begin
                lengths_1 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_2 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h2 == _GEN_182[7:0]) begin
                lengths_2 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_3 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h3 == _GEN_182[7:0]) begin
                lengths_3 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_4 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h4 == _GEN_182[7:0]) begin
                lengths_4 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_5 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h5 == _GEN_182[7:0]) begin
                lengths_5 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_6 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h6 == _GEN_182[7:0]) begin
                lengths_6 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_7 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h7 == _GEN_182[7:0]) begin
                lengths_7 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_8 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h8 == _GEN_182[7:0]) begin
                lengths_8 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_9 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h9 == _GEN_182[7:0]) begin
                lengths_9 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_10 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha == _GEN_182[7:0]) begin
                lengths_10 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_11 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb == _GEN_182[7:0]) begin
                lengths_11 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_12 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc == _GEN_182[7:0]) begin
                lengths_12 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_13 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd == _GEN_182[7:0]) begin
                lengths_13 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_14 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he == _GEN_182[7:0]) begin
                lengths_14 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_15 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf == _GEN_182[7:0]) begin
                lengths_15 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_16 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h10 == _GEN_182[7:0]) begin
                lengths_16 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_17 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h11 == _GEN_182[7:0]) begin
                lengths_17 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_18 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h12 == _GEN_182[7:0]) begin
                lengths_18 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_19 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h13 == _GEN_182[7:0]) begin
                lengths_19 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_20 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h14 == _GEN_182[7:0]) begin
                lengths_20 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_21 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h15 == _GEN_182[7:0]) begin
                lengths_21 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_22 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h16 == _GEN_182[7:0]) begin
                lengths_22 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_23 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h17 == _GEN_182[7:0]) begin
                lengths_23 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_24 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h18 == _GEN_182[7:0]) begin
                lengths_24 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_25 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h19 == _GEN_182[7:0]) begin
                lengths_25 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_26 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h1a == _GEN_182[7:0]) begin
                lengths_26 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_27 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h1b == _GEN_182[7:0]) begin
                lengths_27 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_28 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h1c == _GEN_182[7:0]) begin
                lengths_28 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_29 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h1d == _GEN_182[7:0]) begin
                lengths_29 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_30 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h1e == _GEN_182[7:0]) begin
                lengths_30 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_31 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h1f == _GEN_182[7:0]) begin
                lengths_31 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_32 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h20 == _GEN_182[7:0]) begin
                lengths_32 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_33 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h21 == _GEN_182[7:0]) begin
                lengths_33 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_34 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h22 == _GEN_182[7:0]) begin
                lengths_34 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_35 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h23 == _GEN_182[7:0]) begin
                lengths_35 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_36 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h24 == _GEN_182[7:0]) begin
                lengths_36 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_37 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h25 == _GEN_182[7:0]) begin
                lengths_37 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_38 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h26 == _GEN_182[7:0]) begin
                lengths_38 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_39 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h27 == _GEN_182[7:0]) begin
                lengths_39 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_40 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h28 == _GEN_182[7:0]) begin
                lengths_40 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_41 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h29 == _GEN_182[7:0]) begin
                lengths_41 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_42 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h2a == _GEN_182[7:0]) begin
                lengths_42 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_43 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h2b == _GEN_182[7:0]) begin
                lengths_43 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_44 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h2c == _GEN_182[7:0]) begin
                lengths_44 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_45 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h2d == _GEN_182[7:0]) begin
                lengths_45 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_46 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h2e == _GEN_182[7:0]) begin
                lengths_46 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_47 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h2f == _GEN_182[7:0]) begin
                lengths_47 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_48 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h30 == _GEN_182[7:0]) begin
                lengths_48 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_49 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h31 == _GEN_182[7:0]) begin
                lengths_49 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_50 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h32 == _GEN_182[7:0]) begin
                lengths_50 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_51 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h33 == _GEN_182[7:0]) begin
                lengths_51 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_52 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h34 == _GEN_182[7:0]) begin
                lengths_52 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_53 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h35 == _GEN_182[7:0]) begin
                lengths_53 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_54 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h36 == _GEN_182[7:0]) begin
                lengths_54 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_55 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h37 == _GEN_182[7:0]) begin
                lengths_55 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_56 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h38 == _GEN_182[7:0]) begin
                lengths_56 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_57 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h39 == _GEN_182[7:0]) begin
                lengths_57 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_58 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h3a == _GEN_182[7:0]) begin
                lengths_58 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_59 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h3b == _GEN_182[7:0]) begin
                lengths_59 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_60 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h3c == _GEN_182[7:0]) begin
                lengths_60 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_61 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h3d == _GEN_182[7:0]) begin
                lengths_61 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_62 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h3e == _GEN_182[7:0]) begin
                lengths_62 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_63 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h3f == _GEN_182[7:0]) begin
                lengths_63 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_64 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h40 == _GEN_182[7:0]) begin
                lengths_64 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_65 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h41 == _GEN_182[7:0]) begin
                lengths_65 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_66 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h42 == _GEN_182[7:0]) begin
                lengths_66 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_67 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h43 == _GEN_182[7:0]) begin
                lengths_67 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_68 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h44 == _GEN_182[7:0]) begin
                lengths_68 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_69 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h45 == _GEN_182[7:0]) begin
                lengths_69 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_70 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h46 == _GEN_182[7:0]) begin
                lengths_70 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_71 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h47 == _GEN_182[7:0]) begin
                lengths_71 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_72 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h48 == _GEN_182[7:0]) begin
                lengths_72 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_73 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h49 == _GEN_182[7:0]) begin
                lengths_73 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_74 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h4a == _GEN_182[7:0]) begin
                lengths_74 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_75 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h4b == _GEN_182[7:0]) begin
                lengths_75 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_76 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h4c == _GEN_182[7:0]) begin
                lengths_76 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_77 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h4d == _GEN_182[7:0]) begin
                lengths_77 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_78 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h4e == _GEN_182[7:0]) begin
                lengths_78 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_79 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h4f == _GEN_182[7:0]) begin
                lengths_79 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_80 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h50 == _GEN_182[7:0]) begin
                lengths_80 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_81 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h51 == _GEN_182[7:0]) begin
                lengths_81 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_82 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h52 == _GEN_182[7:0]) begin
                lengths_82 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_83 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h53 == _GEN_182[7:0]) begin
                lengths_83 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_84 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h54 == _GEN_182[7:0]) begin
                lengths_84 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_85 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h55 == _GEN_182[7:0]) begin
                lengths_85 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_86 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h56 == _GEN_182[7:0]) begin
                lengths_86 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_87 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h57 == _GEN_182[7:0]) begin
                lengths_87 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_88 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h58 == _GEN_182[7:0]) begin
                lengths_88 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_89 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h59 == _GEN_182[7:0]) begin
                lengths_89 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_90 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h5a == _GEN_182[7:0]) begin
                lengths_90 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_91 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h5b == _GEN_182[7:0]) begin
                lengths_91 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_92 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h5c == _GEN_182[7:0]) begin
                lengths_92 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_93 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h5d == _GEN_182[7:0]) begin
                lengths_93 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_94 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h5e == _GEN_182[7:0]) begin
                lengths_94 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_95 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h5f == _GEN_182[7:0]) begin
                lengths_95 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_96 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h60 == _GEN_182[7:0]) begin
                lengths_96 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_97 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h61 == _GEN_182[7:0]) begin
                lengths_97 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_98 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h62 == _GEN_182[7:0]) begin
                lengths_98 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_99 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h63 == _GEN_182[7:0]) begin
                lengths_99 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_100 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h64 == _GEN_182[7:0]) begin
                lengths_100 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_101 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h65 == _GEN_182[7:0]) begin
                lengths_101 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_102 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h66 == _GEN_182[7:0]) begin
                lengths_102 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_103 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h67 == _GEN_182[7:0]) begin
                lengths_103 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_104 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h68 == _GEN_182[7:0]) begin
                lengths_104 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_105 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h69 == _GEN_182[7:0]) begin
                lengths_105 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_106 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h6a == _GEN_182[7:0]) begin
                lengths_106 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_107 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h6b == _GEN_182[7:0]) begin
                lengths_107 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_108 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h6c == _GEN_182[7:0]) begin
                lengths_108 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_109 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h6d == _GEN_182[7:0]) begin
                lengths_109 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_110 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h6e == _GEN_182[7:0]) begin
                lengths_110 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_111 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h6f == _GEN_182[7:0]) begin
                lengths_111 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_112 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h70 == _GEN_182[7:0]) begin
                lengths_112 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_113 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h71 == _GEN_182[7:0]) begin
                lengths_113 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_114 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h72 == _GEN_182[7:0]) begin
                lengths_114 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_115 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h73 == _GEN_182[7:0]) begin
                lengths_115 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_116 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h74 == _GEN_182[7:0]) begin
                lengths_116 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_117 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h75 == _GEN_182[7:0]) begin
                lengths_117 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_118 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h76 == _GEN_182[7:0]) begin
                lengths_118 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_119 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h77 == _GEN_182[7:0]) begin
                lengths_119 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_120 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h78 == _GEN_182[7:0]) begin
                lengths_120 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_121 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h79 == _GEN_182[7:0]) begin
                lengths_121 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_122 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h7a == _GEN_182[7:0]) begin
                lengths_122 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_123 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h7b == _GEN_182[7:0]) begin
                lengths_123 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_124 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h7c == _GEN_182[7:0]) begin
                lengths_124 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_125 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h7d == _GEN_182[7:0]) begin
                lengths_125 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_126 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h7e == _GEN_182[7:0]) begin
                lengths_126 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_127 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h7f == _GEN_182[7:0]) begin
                lengths_127 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_128 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h80 == _GEN_182[7:0]) begin
                lengths_128 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_129 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h81 == _GEN_182[7:0]) begin
                lengths_129 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_130 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h82 == _GEN_182[7:0]) begin
                lengths_130 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_131 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h83 == _GEN_182[7:0]) begin
                lengths_131 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_132 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h84 == _GEN_182[7:0]) begin
                lengths_132 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_133 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h85 == _GEN_182[7:0]) begin
                lengths_133 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_134 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h86 == _GEN_182[7:0]) begin
                lengths_134 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_135 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h87 == _GEN_182[7:0]) begin
                lengths_135 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_136 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h88 == _GEN_182[7:0]) begin
                lengths_136 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_137 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h89 == _GEN_182[7:0]) begin
                lengths_137 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_138 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h8a == _GEN_182[7:0]) begin
                lengths_138 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_139 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h8b == _GEN_182[7:0]) begin
                lengths_139 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_140 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h8c == _GEN_182[7:0]) begin
                lengths_140 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_141 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h8d == _GEN_182[7:0]) begin
                lengths_141 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_142 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h8e == _GEN_182[7:0]) begin
                lengths_142 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_143 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h8f == _GEN_182[7:0]) begin
                lengths_143 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_144 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h90 == _GEN_182[7:0]) begin
                lengths_144 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_145 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h91 == _GEN_182[7:0]) begin
                lengths_145 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_146 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h92 == _GEN_182[7:0]) begin
                lengths_146 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_147 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h93 == _GEN_182[7:0]) begin
                lengths_147 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_148 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h94 == _GEN_182[7:0]) begin
                lengths_148 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_149 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h95 == _GEN_182[7:0]) begin
                lengths_149 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_150 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h96 == _GEN_182[7:0]) begin
                lengths_150 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_151 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h97 == _GEN_182[7:0]) begin
                lengths_151 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_152 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h98 == _GEN_182[7:0]) begin
                lengths_152 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_153 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h99 == _GEN_182[7:0]) begin
                lengths_153 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_154 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h9a == _GEN_182[7:0]) begin
                lengths_154 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_155 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h9b == _GEN_182[7:0]) begin
                lengths_155 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_156 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h9c == _GEN_182[7:0]) begin
                lengths_156 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_157 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h9d == _GEN_182[7:0]) begin
                lengths_157 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_158 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h9e == _GEN_182[7:0]) begin
                lengths_158 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_159 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'h9f == _GEN_182[7:0]) begin
                lengths_159 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_160 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha0 == _GEN_182[7:0]) begin
                lengths_160 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_161 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha1 == _GEN_182[7:0]) begin
                lengths_161 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_162 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha2 == _GEN_182[7:0]) begin
                lengths_162 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_163 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha3 == _GEN_182[7:0]) begin
                lengths_163 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_164 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha4 == _GEN_182[7:0]) begin
                lengths_164 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_165 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha5 == _GEN_182[7:0]) begin
                lengths_165 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_166 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha6 == _GEN_182[7:0]) begin
                lengths_166 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_167 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha7 == _GEN_182[7:0]) begin
                lengths_167 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_168 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha8 == _GEN_182[7:0]) begin
                lengths_168 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_169 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'ha9 == _GEN_182[7:0]) begin
                lengths_169 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_170 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'haa == _GEN_182[7:0]) begin
                lengths_170 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_171 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hab == _GEN_182[7:0]) begin
                lengths_171 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_172 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hac == _GEN_182[7:0]) begin
                lengths_172 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_173 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'had == _GEN_182[7:0]) begin
                lengths_173 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_174 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hae == _GEN_182[7:0]) begin
                lengths_174 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_175 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'haf == _GEN_182[7:0]) begin
                lengths_175 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_176 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb0 == _GEN_182[7:0]) begin
                lengths_176 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_177 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb1 == _GEN_182[7:0]) begin
                lengths_177 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_178 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb2 == _GEN_182[7:0]) begin
                lengths_178 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_179 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb3 == _GEN_182[7:0]) begin
                lengths_179 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_180 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb4 == _GEN_182[7:0]) begin
                lengths_180 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_181 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb5 == _GEN_182[7:0]) begin
                lengths_181 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_182 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb6 == _GEN_182[7:0]) begin
                lengths_182 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_183 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb7 == _GEN_182[7:0]) begin
                lengths_183 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_184 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb8 == _GEN_182[7:0]) begin
                lengths_184 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_185 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hb9 == _GEN_182[7:0]) begin
                lengths_185 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_186 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hba == _GEN_182[7:0]) begin
                lengths_186 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_187 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hbb == _GEN_182[7:0]) begin
                lengths_187 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_188 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hbc == _GEN_182[7:0]) begin
                lengths_188 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_189 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hbd == _GEN_182[7:0]) begin
                lengths_189 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_190 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hbe == _GEN_182[7:0]) begin
                lengths_190 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_191 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hbf == _GEN_182[7:0]) begin
                lengths_191 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_192 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc0 == _GEN_182[7:0]) begin
                lengths_192 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_193 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc1 == _GEN_182[7:0]) begin
                lengths_193 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_194 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc2 == _GEN_182[7:0]) begin
                lengths_194 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_195 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc3 == _GEN_182[7:0]) begin
                lengths_195 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_196 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc4 == _GEN_182[7:0]) begin
                lengths_196 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_197 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc5 == _GEN_182[7:0]) begin
                lengths_197 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_198 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc6 == _GEN_182[7:0]) begin
                lengths_198 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_199 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc7 == _GEN_182[7:0]) begin
                lengths_199 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_200 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc8 == _GEN_182[7:0]) begin
                lengths_200 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_201 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hc9 == _GEN_182[7:0]) begin
                lengths_201 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_202 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hca == _GEN_182[7:0]) begin
                lengths_202 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_203 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hcb == _GEN_182[7:0]) begin
                lengths_203 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_204 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hcc == _GEN_182[7:0]) begin
                lengths_204 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_205 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hcd == _GEN_182[7:0]) begin
                lengths_205 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_206 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hce == _GEN_182[7:0]) begin
                lengths_206 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_207 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hcf == _GEN_182[7:0]) begin
                lengths_207 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_208 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd0 == _GEN_182[7:0]) begin
                lengths_208 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_209 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd1 == _GEN_182[7:0]) begin
                lengths_209 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_210 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd2 == _GEN_182[7:0]) begin
                lengths_210 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_211 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd3 == _GEN_182[7:0]) begin
                lengths_211 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_212 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd4 == _GEN_182[7:0]) begin
                lengths_212 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_213 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd5 == _GEN_182[7:0]) begin
                lengths_213 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_214 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd6 == _GEN_182[7:0]) begin
                lengths_214 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_215 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd7 == _GEN_182[7:0]) begin
                lengths_215 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_216 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd8 == _GEN_182[7:0]) begin
                lengths_216 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_217 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hd9 == _GEN_182[7:0]) begin
                lengths_217 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_218 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hda == _GEN_182[7:0]) begin
                lengths_218 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_219 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hdb == _GEN_182[7:0]) begin
                lengths_219 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_220 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hdc == _GEN_182[7:0]) begin
                lengths_220 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_221 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hdd == _GEN_182[7:0]) begin
                lengths_221 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_222 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hde == _GEN_182[7:0]) begin
                lengths_222 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_223 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hdf == _GEN_182[7:0]) begin
                lengths_223 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_224 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he0 == _GEN_182[7:0]) begin
                lengths_224 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_225 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he1 == _GEN_182[7:0]) begin
                lengths_225 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_226 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he2 == _GEN_182[7:0]) begin
                lengths_226 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_227 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he3 == _GEN_182[7:0]) begin
                lengths_227 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_228 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he4 == _GEN_182[7:0]) begin
                lengths_228 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_229 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he5 == _GEN_182[7:0]) begin
                lengths_229 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_230 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he6 == _GEN_182[7:0]) begin
                lengths_230 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_231 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he7 == _GEN_182[7:0]) begin
                lengths_231 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_232 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he8 == _GEN_182[7:0]) begin
                lengths_232 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_233 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'he9 == _GEN_182[7:0]) begin
                lengths_233 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_234 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hea == _GEN_182[7:0]) begin
                lengths_234 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_235 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'heb == _GEN_182[7:0]) begin
                lengths_235 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_236 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hec == _GEN_182[7:0]) begin
                lengths_236 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_237 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hed == _GEN_182[7:0]) begin
                lengths_237 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_238 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hee == _GEN_182[7:0]) begin
                lengths_238 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_239 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hef == _GEN_182[7:0]) begin
                lengths_239 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_240 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf0 == _GEN_182[7:0]) begin
                lengths_240 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_241 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf1 == _GEN_182[7:0]) begin
                lengths_241 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_242 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf2 == _GEN_182[7:0]) begin
                lengths_242 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_243 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf3 == _GEN_182[7:0]) begin
                lengths_243 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_244 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf4 == _GEN_182[7:0]) begin
                lengths_244 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_245 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf5 == _GEN_182[7:0]) begin
                lengths_245 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_246 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf6 == _GEN_182[7:0]) begin
                lengths_246 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_247 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf7 == _GEN_182[7:0]) begin
                lengths_247 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_248 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf8 == _GEN_182[7:0]) begin
                lengths_248 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_249 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hf9 == _GEN_182[7:0]) begin
                lengths_249 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_250 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hfa == _GEN_182[7:0]) begin
                lengths_250 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_251 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hfb == _GEN_182[7:0]) begin
                lengths_251 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_252 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hfc == _GEN_182[7:0]) begin
                lengths_252 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_253 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hfd == _GEN_182[7:0]) begin
                lengths_253 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_254 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hfe == _GEN_182[7:0]) begin
                lengths_254 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      lengths_255 <= 5'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (!(_GEN_182[8])) begin
              if (8'hff == _GEN_182[7:0]) begin
                lengths_255 <= _lengths_T_59;
              end
            end
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h0 == characterIndex) begin
              lengthsOut_0 <= _T_69;
            end
          end else if (8'h0 == characterIndex) begin
            if (8'hff == characterIndex) begin
              lengthsOut_0 <= lengths_255;
            end else if (8'hfe == characterIndex) begin
              lengthsOut_0 <= lengths_254;
            end else if (8'hfd == characterIndex) begin
              lengthsOut_0 <= lengths_253;
            end else if (8'hfc == characterIndex) begin
              lengthsOut_0 <= lengths_252;
            end else if (8'hfb == characterIndex) begin
              lengthsOut_0 <= lengths_251;
            end else if (8'hfa == characterIndex) begin
              lengthsOut_0 <= lengths_250;
            end else if (8'hf9 == characterIndex) begin
              lengthsOut_0 <= lengths_249;
            end else if (8'hf8 == characterIndex) begin
              lengthsOut_0 <= lengths_248;
            end else if (8'hf7 == characterIndex) begin
              lengthsOut_0 <= lengths_247;
            end else if (8'hf6 == characterIndex) begin
              lengthsOut_0 <= lengths_246;
            end else if (8'hf5 == characterIndex) begin
              lengthsOut_0 <= lengths_245;
            end else if (8'hf4 == characterIndex) begin
              lengthsOut_0 <= lengths_244;
            end else if (8'hf3 == characterIndex) begin
              lengthsOut_0 <= lengths_243;
            end else if (8'hf2 == characterIndex) begin
              lengthsOut_0 <= lengths_242;
            end else if (8'hf1 == characterIndex) begin
              lengthsOut_0 <= lengths_241;
            end else if (8'hf0 == characterIndex) begin
              lengthsOut_0 <= lengths_240;
            end else if (8'hef == characterIndex) begin
              lengthsOut_0 <= lengths_239;
            end else if (8'hee == characterIndex) begin
              lengthsOut_0 <= lengths_238;
            end else if (8'hed == characterIndex) begin
              lengthsOut_0 <= lengths_237;
            end else if (8'hec == characterIndex) begin
              lengthsOut_0 <= lengths_236;
            end else if (8'heb == characterIndex) begin
              lengthsOut_0 <= lengths_235;
            end else if (8'hea == characterIndex) begin
              lengthsOut_0 <= lengths_234;
            end else if (8'he9 == characterIndex) begin
              lengthsOut_0 <= lengths_233;
            end else if (8'he8 == characterIndex) begin
              lengthsOut_0 <= lengths_232;
            end else if (8'he7 == characterIndex) begin
              lengthsOut_0 <= lengths_231;
            end else if (8'he6 == characterIndex) begin
              lengthsOut_0 <= lengths_230;
            end else if (8'he5 == characterIndex) begin
              lengthsOut_0 <= lengths_229;
            end else if (8'he4 == characterIndex) begin
              lengthsOut_0 <= lengths_228;
            end else if (8'he3 == characterIndex) begin
              lengthsOut_0 <= lengths_227;
            end else if (8'he2 == characterIndex) begin
              lengthsOut_0 <= lengths_226;
            end else if (8'he1 == characterIndex) begin
              lengthsOut_0 <= lengths_225;
            end else if (8'he0 == characterIndex) begin
              lengthsOut_0 <= lengths_224;
            end else if (8'hdf == characterIndex) begin
              lengthsOut_0 <= lengths_223;
            end else if (8'hde == characterIndex) begin
              lengthsOut_0 <= lengths_222;
            end else if (8'hdd == characterIndex) begin
              lengthsOut_0 <= lengths_221;
            end else if (8'hdc == characterIndex) begin
              lengthsOut_0 <= lengths_220;
            end else if (8'hdb == characterIndex) begin
              lengthsOut_0 <= lengths_219;
            end else if (8'hda == characterIndex) begin
              lengthsOut_0 <= lengths_218;
            end else if (8'hd9 == characterIndex) begin
              lengthsOut_0 <= lengths_217;
            end else if (8'hd8 == characterIndex) begin
              lengthsOut_0 <= lengths_216;
            end else if (8'hd7 == characterIndex) begin
              lengthsOut_0 <= lengths_215;
            end else if (8'hd6 == characterIndex) begin
              lengthsOut_0 <= lengths_214;
            end else if (8'hd5 == characterIndex) begin
              lengthsOut_0 <= lengths_213;
            end else if (8'hd4 == characterIndex) begin
              lengthsOut_0 <= lengths_212;
            end else if (8'hd3 == characterIndex) begin
              lengthsOut_0 <= lengths_211;
            end else if (8'hd2 == characterIndex) begin
              lengthsOut_0 <= lengths_210;
            end else if (8'hd1 == characterIndex) begin
              lengthsOut_0 <= lengths_209;
            end else if (8'hd0 == characterIndex) begin
              lengthsOut_0 <= lengths_208;
            end else if (8'hcf == characterIndex) begin
              lengthsOut_0 <= lengths_207;
            end else if (8'hce == characterIndex) begin
              lengthsOut_0 <= lengths_206;
            end else if (8'hcd == characterIndex) begin
              lengthsOut_0 <= lengths_205;
            end else if (8'hcc == characterIndex) begin
              lengthsOut_0 <= lengths_204;
            end else if (8'hcb == characterIndex) begin
              lengthsOut_0 <= lengths_203;
            end else if (8'hca == characterIndex) begin
              lengthsOut_0 <= lengths_202;
            end else if (8'hc9 == characterIndex) begin
              lengthsOut_0 <= lengths_201;
            end else if (8'hc8 == characterIndex) begin
              lengthsOut_0 <= lengths_200;
            end else if (8'hc7 == characterIndex) begin
              lengthsOut_0 <= lengths_199;
            end else if (8'hc6 == characterIndex) begin
              lengthsOut_0 <= lengths_198;
            end else if (8'hc5 == characterIndex) begin
              lengthsOut_0 <= lengths_197;
            end else if (8'hc4 == characterIndex) begin
              lengthsOut_0 <= lengths_196;
            end else if (8'hc3 == characterIndex) begin
              lengthsOut_0 <= lengths_195;
            end else if (8'hc2 == characterIndex) begin
              lengthsOut_0 <= lengths_194;
            end else if (8'hc1 == characterIndex) begin
              lengthsOut_0 <= lengths_193;
            end else if (8'hc0 == characterIndex) begin
              lengthsOut_0 <= lengths_192;
            end else if (8'hbf == characterIndex) begin
              lengthsOut_0 <= lengths_191;
            end else if (8'hbe == characterIndex) begin
              lengthsOut_0 <= lengths_190;
            end else if (8'hbd == characterIndex) begin
              lengthsOut_0 <= lengths_189;
            end else if (8'hbc == characterIndex) begin
              lengthsOut_0 <= lengths_188;
            end else if (8'hbb == characterIndex) begin
              lengthsOut_0 <= lengths_187;
            end else if (8'hba == characterIndex) begin
              lengthsOut_0 <= lengths_186;
            end else if (8'hb9 == characterIndex) begin
              lengthsOut_0 <= lengths_185;
            end else if (8'hb8 == characterIndex) begin
              lengthsOut_0 <= lengths_184;
            end else if (8'hb7 == characterIndex) begin
              lengthsOut_0 <= lengths_183;
            end else if (8'hb6 == characterIndex) begin
              lengthsOut_0 <= lengths_182;
            end else if (8'hb5 == characterIndex) begin
              lengthsOut_0 <= lengths_181;
            end else if (8'hb4 == characterIndex) begin
              lengthsOut_0 <= lengths_180;
            end else if (8'hb3 == characterIndex) begin
              lengthsOut_0 <= lengths_179;
            end else if (8'hb2 == characterIndex) begin
              lengthsOut_0 <= lengths_178;
            end else if (8'hb1 == characterIndex) begin
              lengthsOut_0 <= lengths_177;
            end else if (8'hb0 == characterIndex) begin
              lengthsOut_0 <= lengths_176;
            end else if (8'haf == characterIndex) begin
              lengthsOut_0 <= lengths_175;
            end else if (8'hae == characterIndex) begin
              lengthsOut_0 <= lengths_174;
            end else if (8'had == characterIndex) begin
              lengthsOut_0 <= lengths_173;
            end else if (8'hac == characterIndex) begin
              lengthsOut_0 <= lengths_172;
            end else if (8'hab == characterIndex) begin
              lengthsOut_0 <= lengths_171;
            end else if (8'haa == characterIndex) begin
              lengthsOut_0 <= lengths_170;
            end else if (8'ha9 == characterIndex) begin
              lengthsOut_0 <= lengths_169;
            end else if (8'ha8 == characterIndex) begin
              lengthsOut_0 <= lengths_168;
            end else if (8'ha7 == characterIndex) begin
              lengthsOut_0 <= lengths_167;
            end else if (8'ha6 == characterIndex) begin
              lengthsOut_0 <= lengths_166;
            end else if (8'ha5 == characterIndex) begin
              lengthsOut_0 <= lengths_165;
            end else if (8'ha4 == characterIndex) begin
              lengthsOut_0 <= lengths_164;
            end else if (8'ha3 == characterIndex) begin
              lengthsOut_0 <= lengths_163;
            end else if (8'ha2 == characterIndex) begin
              lengthsOut_0 <= lengths_162;
            end else if (8'ha1 == characterIndex) begin
              lengthsOut_0 <= lengths_161;
            end else if (8'ha0 == characterIndex) begin
              lengthsOut_0 <= lengths_160;
            end else if (8'h9f == characterIndex) begin
              lengthsOut_0 <= lengths_159;
            end else if (8'h9e == characterIndex) begin
              lengthsOut_0 <= lengths_158;
            end else if (8'h9d == characterIndex) begin
              lengthsOut_0 <= lengths_157;
            end else if (8'h9c == characterIndex) begin
              lengthsOut_0 <= lengths_156;
            end else if (8'h9b == characterIndex) begin
              lengthsOut_0 <= lengths_155;
            end else if (8'h9a == characterIndex) begin
              lengthsOut_0 <= lengths_154;
            end else if (8'h99 == characterIndex) begin
              lengthsOut_0 <= lengths_153;
            end else if (8'h98 == characterIndex) begin
              lengthsOut_0 <= lengths_152;
            end else if (8'h97 == characterIndex) begin
              lengthsOut_0 <= lengths_151;
            end else if (8'h96 == characterIndex) begin
              lengthsOut_0 <= lengths_150;
            end else if (8'h95 == characterIndex) begin
              lengthsOut_0 <= lengths_149;
            end else if (8'h94 == characterIndex) begin
              lengthsOut_0 <= lengths_148;
            end else if (8'h93 == characterIndex) begin
              lengthsOut_0 <= lengths_147;
            end else if (8'h92 == characterIndex) begin
              lengthsOut_0 <= lengths_146;
            end else if (8'h91 == characterIndex) begin
              lengthsOut_0 <= lengths_145;
            end else if (8'h90 == characterIndex) begin
              lengthsOut_0 <= lengths_144;
            end else if (8'h8f == characterIndex) begin
              lengthsOut_0 <= lengths_143;
            end else if (8'h8e == characterIndex) begin
              lengthsOut_0 <= lengths_142;
            end else if (8'h8d == characterIndex) begin
              lengthsOut_0 <= lengths_141;
            end else if (8'h8c == characterIndex) begin
              lengthsOut_0 <= lengths_140;
            end else if (8'h8b == characterIndex) begin
              lengthsOut_0 <= lengths_139;
            end else if (8'h8a == characterIndex) begin
              lengthsOut_0 <= lengths_138;
            end else if (8'h89 == characterIndex) begin
              lengthsOut_0 <= lengths_137;
            end else if (8'h88 == characterIndex) begin
              lengthsOut_0 <= lengths_136;
            end else if (8'h87 == characterIndex) begin
              lengthsOut_0 <= lengths_135;
            end else if (8'h86 == characterIndex) begin
              lengthsOut_0 <= lengths_134;
            end else if (8'h85 == characterIndex) begin
              lengthsOut_0 <= lengths_133;
            end else if (8'h84 == characterIndex) begin
              lengthsOut_0 <= lengths_132;
            end else if (8'h83 == characterIndex) begin
              lengthsOut_0 <= lengths_131;
            end else if (8'h82 == characterIndex) begin
              lengthsOut_0 <= lengths_130;
            end else if (8'h81 == characterIndex) begin
              lengthsOut_0 <= lengths_129;
            end else if (8'h80 == characterIndex) begin
              lengthsOut_0 <= lengths_128;
            end else if (8'h7f == characterIndex) begin
              lengthsOut_0 <= lengths_127;
            end else if (8'h7e == characterIndex) begin
              lengthsOut_0 <= lengths_126;
            end else if (8'h7d == characterIndex) begin
              lengthsOut_0 <= lengths_125;
            end else if (8'h7c == characterIndex) begin
              lengthsOut_0 <= lengths_124;
            end else if (8'h7b == characterIndex) begin
              lengthsOut_0 <= lengths_123;
            end else if (8'h7a == characterIndex) begin
              lengthsOut_0 <= lengths_122;
            end else if (8'h79 == characterIndex) begin
              lengthsOut_0 <= lengths_121;
            end else if (8'h78 == characterIndex) begin
              lengthsOut_0 <= lengths_120;
            end else if (8'h77 == characterIndex) begin
              lengthsOut_0 <= lengths_119;
            end else if (8'h76 == characterIndex) begin
              lengthsOut_0 <= lengths_118;
            end else if (8'h75 == characterIndex) begin
              lengthsOut_0 <= lengths_117;
            end else if (8'h74 == characterIndex) begin
              lengthsOut_0 <= lengths_116;
            end else if (8'h73 == characterIndex) begin
              lengthsOut_0 <= lengths_115;
            end else if (8'h72 == characterIndex) begin
              lengthsOut_0 <= lengths_114;
            end else if (8'h71 == characterIndex) begin
              lengthsOut_0 <= lengths_113;
            end else if (8'h70 == characterIndex) begin
              lengthsOut_0 <= lengths_112;
            end else if (8'h6f == characterIndex) begin
              lengthsOut_0 <= lengths_111;
            end else if (8'h6e == characterIndex) begin
              lengthsOut_0 <= lengths_110;
            end else if (8'h6d == characterIndex) begin
              lengthsOut_0 <= lengths_109;
            end else if (8'h6c == characterIndex) begin
              lengthsOut_0 <= lengths_108;
            end else if (8'h6b == characterIndex) begin
              lengthsOut_0 <= lengths_107;
            end else if (8'h6a == characterIndex) begin
              lengthsOut_0 <= lengths_106;
            end else if (8'h69 == characterIndex) begin
              lengthsOut_0 <= lengths_105;
            end else if (8'h68 == characterIndex) begin
              lengthsOut_0 <= lengths_104;
            end else if (8'h67 == characterIndex) begin
              lengthsOut_0 <= lengths_103;
            end else if (8'h66 == characterIndex) begin
              lengthsOut_0 <= lengths_102;
            end else if (8'h65 == characterIndex) begin
              lengthsOut_0 <= lengths_101;
            end else if (8'h64 == characterIndex) begin
              lengthsOut_0 <= lengths_100;
            end else if (8'h63 == characterIndex) begin
              lengthsOut_0 <= lengths_99;
            end else if (8'h62 == characterIndex) begin
              lengthsOut_0 <= lengths_98;
            end else if (8'h61 == characterIndex) begin
              lengthsOut_0 <= lengths_97;
            end else if (8'h60 == characterIndex) begin
              lengthsOut_0 <= lengths_96;
            end else if (8'h5f == characterIndex) begin
              lengthsOut_0 <= lengths_95;
            end else if (8'h5e == characterIndex) begin
              lengthsOut_0 <= lengths_94;
            end else if (8'h5d == characterIndex) begin
              lengthsOut_0 <= lengths_93;
            end else if (8'h5c == characterIndex) begin
              lengthsOut_0 <= lengths_92;
            end else if (8'h5b == characterIndex) begin
              lengthsOut_0 <= lengths_91;
            end else if (8'h5a == characterIndex) begin
              lengthsOut_0 <= lengths_90;
            end else if (8'h59 == characterIndex) begin
              lengthsOut_0 <= lengths_89;
            end else if (8'h58 == characterIndex) begin
              lengthsOut_0 <= lengths_88;
            end else if (8'h57 == characterIndex) begin
              lengthsOut_0 <= lengths_87;
            end else if (8'h56 == characterIndex) begin
              lengthsOut_0 <= lengths_86;
            end else if (8'h55 == characterIndex) begin
              lengthsOut_0 <= lengths_85;
            end else if (8'h54 == characterIndex) begin
              lengthsOut_0 <= lengths_84;
            end else if (8'h53 == characterIndex) begin
              lengthsOut_0 <= lengths_83;
            end else if (8'h52 == characterIndex) begin
              lengthsOut_0 <= lengths_82;
            end else if (8'h51 == characterIndex) begin
              lengthsOut_0 <= lengths_81;
            end else if (8'h50 == characterIndex) begin
              lengthsOut_0 <= lengths_80;
            end else if (8'h4f == characterIndex) begin
              lengthsOut_0 <= lengths_79;
            end else if (8'h4e == characterIndex) begin
              lengthsOut_0 <= lengths_78;
            end else if (8'h4d == characterIndex) begin
              lengthsOut_0 <= lengths_77;
            end else if (8'h4c == characterIndex) begin
              lengthsOut_0 <= lengths_76;
            end else if (8'h4b == characterIndex) begin
              lengthsOut_0 <= lengths_75;
            end else if (8'h4a == characterIndex) begin
              lengthsOut_0 <= lengths_74;
            end else if (8'h49 == characterIndex) begin
              lengthsOut_0 <= lengths_73;
            end else if (8'h48 == characterIndex) begin
              lengthsOut_0 <= lengths_72;
            end else if (8'h47 == characterIndex) begin
              lengthsOut_0 <= lengths_71;
            end else if (8'h46 == characterIndex) begin
              lengthsOut_0 <= lengths_70;
            end else if (8'h45 == characterIndex) begin
              lengthsOut_0 <= lengths_69;
            end else if (8'h44 == characterIndex) begin
              lengthsOut_0 <= lengths_68;
            end else if (8'h43 == characterIndex) begin
              lengthsOut_0 <= lengths_67;
            end else if (8'h42 == characterIndex) begin
              lengthsOut_0 <= lengths_66;
            end else if (8'h41 == characterIndex) begin
              lengthsOut_0 <= lengths_65;
            end else if (8'h40 == characterIndex) begin
              lengthsOut_0 <= lengths_64;
            end else if (8'h3f == characterIndex) begin
              lengthsOut_0 <= lengths_63;
            end else if (8'h3e == characterIndex) begin
              lengthsOut_0 <= lengths_62;
            end else if (8'h3d == characterIndex) begin
              lengthsOut_0 <= lengths_61;
            end else if (8'h3c == characterIndex) begin
              lengthsOut_0 <= lengths_60;
            end else if (8'h3b == characterIndex) begin
              lengthsOut_0 <= lengths_59;
            end else if (8'h3a == characterIndex) begin
              lengthsOut_0 <= lengths_58;
            end else if (8'h39 == characterIndex) begin
              lengthsOut_0 <= lengths_57;
            end else if (8'h38 == characterIndex) begin
              lengthsOut_0 <= lengths_56;
            end else if (8'h37 == characterIndex) begin
              lengthsOut_0 <= lengths_55;
            end else if (8'h36 == characterIndex) begin
              lengthsOut_0 <= lengths_54;
            end else if (8'h35 == characterIndex) begin
              lengthsOut_0 <= lengths_53;
            end else if (8'h34 == characterIndex) begin
              lengthsOut_0 <= lengths_52;
            end else if (8'h33 == characterIndex) begin
              lengthsOut_0 <= lengths_51;
            end else if (8'h32 == characterIndex) begin
              lengthsOut_0 <= lengths_50;
            end else if (8'h31 == characterIndex) begin
              lengthsOut_0 <= lengths_49;
            end else if (8'h30 == characterIndex) begin
              lengthsOut_0 <= lengths_48;
            end else if (8'h2f == characterIndex) begin
              lengthsOut_0 <= lengths_47;
            end else if (8'h2e == characterIndex) begin
              lengthsOut_0 <= lengths_46;
            end else if (8'h2d == characterIndex) begin
              lengthsOut_0 <= lengths_45;
            end else if (8'h2c == characterIndex) begin
              lengthsOut_0 <= lengths_44;
            end else if (8'h2b == characterIndex) begin
              lengthsOut_0 <= lengths_43;
            end else if (8'h2a == characterIndex) begin
              lengthsOut_0 <= lengths_42;
            end else if (8'h29 == characterIndex) begin
              lengthsOut_0 <= lengths_41;
            end else if (8'h28 == characterIndex) begin
              lengthsOut_0 <= lengths_40;
            end else if (8'h27 == characterIndex) begin
              lengthsOut_0 <= lengths_39;
            end else if (8'h26 == characterIndex) begin
              lengthsOut_0 <= lengths_38;
            end else if (8'h25 == characterIndex) begin
              lengthsOut_0 <= lengths_37;
            end else if (8'h24 == characterIndex) begin
              lengthsOut_0 <= lengths_36;
            end else if (8'h23 == characterIndex) begin
              lengthsOut_0 <= lengths_35;
            end else if (8'h22 == characterIndex) begin
              lengthsOut_0 <= lengths_34;
            end else if (8'h21 == characterIndex) begin
              lengthsOut_0 <= lengths_33;
            end else if (8'h20 == characterIndex) begin
              lengthsOut_0 <= lengths_32;
            end else if (8'h1f == characterIndex) begin
              lengthsOut_0 <= lengths_31;
            end else if (8'h1e == characterIndex) begin
              lengthsOut_0 <= lengths_30;
            end else if (8'h1d == characterIndex) begin
              lengthsOut_0 <= lengths_29;
            end else if (8'h1c == characterIndex) begin
              lengthsOut_0 <= lengths_28;
            end else if (8'h1b == characterIndex) begin
              lengthsOut_0 <= lengths_27;
            end else if (8'h1a == characterIndex) begin
              lengthsOut_0 <= lengths_26;
            end else if (8'h19 == characterIndex) begin
              lengthsOut_0 <= lengths_25;
            end else if (8'h18 == characterIndex) begin
              lengthsOut_0 <= lengths_24;
            end else if (8'h17 == characterIndex) begin
              lengthsOut_0 <= lengths_23;
            end else if (8'h16 == characterIndex) begin
              lengthsOut_0 <= lengths_22;
            end else if (8'h15 == characterIndex) begin
              lengthsOut_0 <= lengths_21;
            end else if (8'h14 == characterIndex) begin
              lengthsOut_0 <= lengths_20;
            end else if (8'h13 == characterIndex) begin
              lengthsOut_0 <= lengths_19;
            end else if (8'h12 == characterIndex) begin
              lengthsOut_0 <= lengths_18;
            end else if (8'h11 == characterIndex) begin
              lengthsOut_0 <= lengths_17;
            end else if (8'h10 == characterIndex) begin
              lengthsOut_0 <= lengths_16;
            end else if (8'hf == characterIndex) begin
              lengthsOut_0 <= lengths_15;
            end else if (8'he == characterIndex) begin
              lengthsOut_0 <= lengths_14;
            end else if (8'hd == characterIndex) begin
              lengthsOut_0 <= lengths_13;
            end else if (8'hc == characterIndex) begin
              lengthsOut_0 <= lengths_12;
            end else if (8'hb == characterIndex) begin
              lengthsOut_0 <= lengths_11;
            end else if (8'ha == characterIndex) begin
              lengthsOut_0 <= lengths_10;
            end else if (8'h9 == characterIndex) begin
              lengthsOut_0 <= lengths_9;
            end else if (8'h8 == characterIndex) begin
              lengthsOut_0 <= lengths_8;
            end else if (8'h7 == characterIndex) begin
              lengthsOut_0 <= lengths_7;
            end else if (8'h6 == characterIndex) begin
              lengthsOut_0 <= lengths_6;
            end else if (8'h5 == characterIndex) begin
              lengthsOut_0 <= lengths_5;
            end else if (8'h4 == characterIndex) begin
              lengthsOut_0 <= lengths_4;
            end else if (8'h3 == characterIndex) begin
              lengthsOut_0 <= lengths_3;
            end else if (8'h2 == characterIndex) begin
              lengthsOut_0 <= lengths_2;
            end else if (8'h1 == characterIndex) begin
              lengthsOut_0 <= lengths_1;
            end else begin
              lengthsOut_0 <= lengths_0;
            end
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h1 == characterIndex) begin
              lengthsOut_1 <= _T_69;
            end
          end else if (8'h1 == characterIndex) begin
            if (8'hff == characterIndex) begin
              lengthsOut_1 <= lengths_255;
            end else if (8'hfe == characterIndex) begin
              lengthsOut_1 <= lengths_254;
            end else if (8'hfd == characterIndex) begin
              lengthsOut_1 <= lengths_253;
            end else if (8'hfc == characterIndex) begin
              lengthsOut_1 <= lengths_252;
            end else if (8'hfb == characterIndex) begin
              lengthsOut_1 <= lengths_251;
            end else if (8'hfa == characterIndex) begin
              lengthsOut_1 <= lengths_250;
            end else if (8'hf9 == characterIndex) begin
              lengthsOut_1 <= lengths_249;
            end else if (8'hf8 == characterIndex) begin
              lengthsOut_1 <= lengths_248;
            end else if (8'hf7 == characterIndex) begin
              lengthsOut_1 <= lengths_247;
            end else if (8'hf6 == characterIndex) begin
              lengthsOut_1 <= lengths_246;
            end else if (8'hf5 == characterIndex) begin
              lengthsOut_1 <= lengths_245;
            end else if (8'hf4 == characterIndex) begin
              lengthsOut_1 <= lengths_244;
            end else if (8'hf3 == characterIndex) begin
              lengthsOut_1 <= lengths_243;
            end else if (8'hf2 == characterIndex) begin
              lengthsOut_1 <= lengths_242;
            end else if (8'hf1 == characterIndex) begin
              lengthsOut_1 <= lengths_241;
            end else if (8'hf0 == characterIndex) begin
              lengthsOut_1 <= lengths_240;
            end else if (8'hef == characterIndex) begin
              lengthsOut_1 <= lengths_239;
            end else if (8'hee == characterIndex) begin
              lengthsOut_1 <= lengths_238;
            end else if (8'hed == characterIndex) begin
              lengthsOut_1 <= lengths_237;
            end else if (8'hec == characterIndex) begin
              lengthsOut_1 <= lengths_236;
            end else if (8'heb == characterIndex) begin
              lengthsOut_1 <= lengths_235;
            end else if (8'hea == characterIndex) begin
              lengthsOut_1 <= lengths_234;
            end else if (8'he9 == characterIndex) begin
              lengthsOut_1 <= lengths_233;
            end else if (8'he8 == characterIndex) begin
              lengthsOut_1 <= lengths_232;
            end else if (8'he7 == characterIndex) begin
              lengthsOut_1 <= lengths_231;
            end else if (8'he6 == characterIndex) begin
              lengthsOut_1 <= lengths_230;
            end else if (8'he5 == characterIndex) begin
              lengthsOut_1 <= lengths_229;
            end else if (8'he4 == characterIndex) begin
              lengthsOut_1 <= lengths_228;
            end else if (8'he3 == characterIndex) begin
              lengthsOut_1 <= lengths_227;
            end else if (8'he2 == characterIndex) begin
              lengthsOut_1 <= lengths_226;
            end else if (8'he1 == characterIndex) begin
              lengthsOut_1 <= lengths_225;
            end else if (8'he0 == characterIndex) begin
              lengthsOut_1 <= lengths_224;
            end else if (8'hdf == characterIndex) begin
              lengthsOut_1 <= lengths_223;
            end else if (8'hde == characterIndex) begin
              lengthsOut_1 <= lengths_222;
            end else if (8'hdd == characterIndex) begin
              lengthsOut_1 <= lengths_221;
            end else if (8'hdc == characterIndex) begin
              lengthsOut_1 <= lengths_220;
            end else if (8'hdb == characterIndex) begin
              lengthsOut_1 <= lengths_219;
            end else if (8'hda == characterIndex) begin
              lengthsOut_1 <= lengths_218;
            end else if (8'hd9 == characterIndex) begin
              lengthsOut_1 <= lengths_217;
            end else if (8'hd8 == characterIndex) begin
              lengthsOut_1 <= lengths_216;
            end else if (8'hd7 == characterIndex) begin
              lengthsOut_1 <= lengths_215;
            end else if (8'hd6 == characterIndex) begin
              lengthsOut_1 <= lengths_214;
            end else if (8'hd5 == characterIndex) begin
              lengthsOut_1 <= lengths_213;
            end else if (8'hd4 == characterIndex) begin
              lengthsOut_1 <= lengths_212;
            end else if (8'hd3 == characterIndex) begin
              lengthsOut_1 <= lengths_211;
            end else if (8'hd2 == characterIndex) begin
              lengthsOut_1 <= lengths_210;
            end else if (8'hd1 == characterIndex) begin
              lengthsOut_1 <= lengths_209;
            end else if (8'hd0 == characterIndex) begin
              lengthsOut_1 <= lengths_208;
            end else if (8'hcf == characterIndex) begin
              lengthsOut_1 <= lengths_207;
            end else if (8'hce == characterIndex) begin
              lengthsOut_1 <= lengths_206;
            end else if (8'hcd == characterIndex) begin
              lengthsOut_1 <= lengths_205;
            end else if (8'hcc == characterIndex) begin
              lengthsOut_1 <= lengths_204;
            end else if (8'hcb == characterIndex) begin
              lengthsOut_1 <= lengths_203;
            end else if (8'hca == characterIndex) begin
              lengthsOut_1 <= lengths_202;
            end else if (8'hc9 == characterIndex) begin
              lengthsOut_1 <= lengths_201;
            end else if (8'hc8 == characterIndex) begin
              lengthsOut_1 <= lengths_200;
            end else if (8'hc7 == characterIndex) begin
              lengthsOut_1 <= lengths_199;
            end else if (8'hc6 == characterIndex) begin
              lengthsOut_1 <= lengths_198;
            end else if (8'hc5 == characterIndex) begin
              lengthsOut_1 <= lengths_197;
            end else if (8'hc4 == characterIndex) begin
              lengthsOut_1 <= lengths_196;
            end else if (8'hc3 == characterIndex) begin
              lengthsOut_1 <= lengths_195;
            end else if (8'hc2 == characterIndex) begin
              lengthsOut_1 <= lengths_194;
            end else if (8'hc1 == characterIndex) begin
              lengthsOut_1 <= lengths_193;
            end else if (8'hc0 == characterIndex) begin
              lengthsOut_1 <= lengths_192;
            end else if (8'hbf == characterIndex) begin
              lengthsOut_1 <= lengths_191;
            end else if (8'hbe == characterIndex) begin
              lengthsOut_1 <= lengths_190;
            end else if (8'hbd == characterIndex) begin
              lengthsOut_1 <= lengths_189;
            end else if (8'hbc == characterIndex) begin
              lengthsOut_1 <= lengths_188;
            end else if (8'hbb == characterIndex) begin
              lengthsOut_1 <= lengths_187;
            end else if (8'hba == characterIndex) begin
              lengthsOut_1 <= lengths_186;
            end else if (8'hb9 == characterIndex) begin
              lengthsOut_1 <= lengths_185;
            end else if (8'hb8 == characterIndex) begin
              lengthsOut_1 <= lengths_184;
            end else if (8'hb7 == characterIndex) begin
              lengthsOut_1 <= lengths_183;
            end else if (8'hb6 == characterIndex) begin
              lengthsOut_1 <= lengths_182;
            end else if (8'hb5 == characterIndex) begin
              lengthsOut_1 <= lengths_181;
            end else if (8'hb4 == characterIndex) begin
              lengthsOut_1 <= lengths_180;
            end else if (8'hb3 == characterIndex) begin
              lengthsOut_1 <= lengths_179;
            end else if (8'hb2 == characterIndex) begin
              lengthsOut_1 <= lengths_178;
            end else if (8'hb1 == characterIndex) begin
              lengthsOut_1 <= lengths_177;
            end else if (8'hb0 == characterIndex) begin
              lengthsOut_1 <= lengths_176;
            end else if (8'haf == characterIndex) begin
              lengthsOut_1 <= lengths_175;
            end else if (8'hae == characterIndex) begin
              lengthsOut_1 <= lengths_174;
            end else if (8'had == characterIndex) begin
              lengthsOut_1 <= lengths_173;
            end else if (8'hac == characterIndex) begin
              lengthsOut_1 <= lengths_172;
            end else if (8'hab == characterIndex) begin
              lengthsOut_1 <= lengths_171;
            end else if (8'haa == characterIndex) begin
              lengthsOut_1 <= lengths_170;
            end else if (8'ha9 == characterIndex) begin
              lengthsOut_1 <= lengths_169;
            end else if (8'ha8 == characterIndex) begin
              lengthsOut_1 <= lengths_168;
            end else if (8'ha7 == characterIndex) begin
              lengthsOut_1 <= lengths_167;
            end else if (8'ha6 == characterIndex) begin
              lengthsOut_1 <= lengths_166;
            end else if (8'ha5 == characterIndex) begin
              lengthsOut_1 <= lengths_165;
            end else if (8'ha4 == characterIndex) begin
              lengthsOut_1 <= lengths_164;
            end else if (8'ha3 == characterIndex) begin
              lengthsOut_1 <= lengths_163;
            end else if (8'ha2 == characterIndex) begin
              lengthsOut_1 <= lengths_162;
            end else if (8'ha1 == characterIndex) begin
              lengthsOut_1 <= lengths_161;
            end else if (8'ha0 == characterIndex) begin
              lengthsOut_1 <= lengths_160;
            end else if (8'h9f == characterIndex) begin
              lengthsOut_1 <= lengths_159;
            end else if (8'h9e == characterIndex) begin
              lengthsOut_1 <= lengths_158;
            end else if (8'h9d == characterIndex) begin
              lengthsOut_1 <= lengths_157;
            end else if (8'h9c == characterIndex) begin
              lengthsOut_1 <= lengths_156;
            end else if (8'h9b == characterIndex) begin
              lengthsOut_1 <= lengths_155;
            end else if (8'h9a == characterIndex) begin
              lengthsOut_1 <= lengths_154;
            end else if (8'h99 == characterIndex) begin
              lengthsOut_1 <= lengths_153;
            end else if (8'h98 == characterIndex) begin
              lengthsOut_1 <= lengths_152;
            end else if (8'h97 == characterIndex) begin
              lengthsOut_1 <= lengths_151;
            end else if (8'h96 == characterIndex) begin
              lengthsOut_1 <= lengths_150;
            end else if (8'h95 == characterIndex) begin
              lengthsOut_1 <= lengths_149;
            end else if (8'h94 == characterIndex) begin
              lengthsOut_1 <= lengths_148;
            end else if (8'h93 == characterIndex) begin
              lengthsOut_1 <= lengths_147;
            end else if (8'h92 == characterIndex) begin
              lengthsOut_1 <= lengths_146;
            end else if (8'h91 == characterIndex) begin
              lengthsOut_1 <= lengths_145;
            end else if (8'h90 == characterIndex) begin
              lengthsOut_1 <= lengths_144;
            end else if (8'h8f == characterIndex) begin
              lengthsOut_1 <= lengths_143;
            end else if (8'h8e == characterIndex) begin
              lengthsOut_1 <= lengths_142;
            end else if (8'h8d == characterIndex) begin
              lengthsOut_1 <= lengths_141;
            end else if (8'h8c == characterIndex) begin
              lengthsOut_1 <= lengths_140;
            end else if (8'h8b == characterIndex) begin
              lengthsOut_1 <= lengths_139;
            end else if (8'h8a == characterIndex) begin
              lengthsOut_1 <= lengths_138;
            end else if (8'h89 == characterIndex) begin
              lengthsOut_1 <= lengths_137;
            end else if (8'h88 == characterIndex) begin
              lengthsOut_1 <= lengths_136;
            end else if (8'h87 == characterIndex) begin
              lengthsOut_1 <= lengths_135;
            end else if (8'h86 == characterIndex) begin
              lengthsOut_1 <= lengths_134;
            end else if (8'h85 == characterIndex) begin
              lengthsOut_1 <= lengths_133;
            end else if (8'h84 == characterIndex) begin
              lengthsOut_1 <= lengths_132;
            end else if (8'h83 == characterIndex) begin
              lengthsOut_1 <= lengths_131;
            end else if (8'h82 == characterIndex) begin
              lengthsOut_1 <= lengths_130;
            end else if (8'h81 == characterIndex) begin
              lengthsOut_1 <= lengths_129;
            end else if (8'h80 == characterIndex) begin
              lengthsOut_1 <= lengths_128;
            end else if (8'h7f == characterIndex) begin
              lengthsOut_1 <= lengths_127;
            end else if (8'h7e == characterIndex) begin
              lengthsOut_1 <= lengths_126;
            end else if (8'h7d == characterIndex) begin
              lengthsOut_1 <= lengths_125;
            end else if (8'h7c == characterIndex) begin
              lengthsOut_1 <= lengths_124;
            end else if (8'h7b == characterIndex) begin
              lengthsOut_1 <= lengths_123;
            end else if (8'h7a == characterIndex) begin
              lengthsOut_1 <= lengths_122;
            end else if (8'h79 == characterIndex) begin
              lengthsOut_1 <= lengths_121;
            end else if (8'h78 == characterIndex) begin
              lengthsOut_1 <= lengths_120;
            end else if (8'h77 == characterIndex) begin
              lengthsOut_1 <= lengths_119;
            end else if (8'h76 == characterIndex) begin
              lengthsOut_1 <= lengths_118;
            end else if (8'h75 == characterIndex) begin
              lengthsOut_1 <= lengths_117;
            end else if (8'h74 == characterIndex) begin
              lengthsOut_1 <= lengths_116;
            end else if (8'h73 == characterIndex) begin
              lengthsOut_1 <= lengths_115;
            end else if (8'h72 == characterIndex) begin
              lengthsOut_1 <= lengths_114;
            end else if (8'h71 == characterIndex) begin
              lengthsOut_1 <= lengths_113;
            end else if (8'h70 == characterIndex) begin
              lengthsOut_1 <= lengths_112;
            end else if (8'h6f == characterIndex) begin
              lengthsOut_1 <= lengths_111;
            end else if (8'h6e == characterIndex) begin
              lengthsOut_1 <= lengths_110;
            end else if (8'h6d == characterIndex) begin
              lengthsOut_1 <= lengths_109;
            end else if (8'h6c == characterIndex) begin
              lengthsOut_1 <= lengths_108;
            end else if (8'h6b == characterIndex) begin
              lengthsOut_1 <= lengths_107;
            end else if (8'h6a == characterIndex) begin
              lengthsOut_1 <= lengths_106;
            end else if (8'h69 == characterIndex) begin
              lengthsOut_1 <= lengths_105;
            end else if (8'h68 == characterIndex) begin
              lengthsOut_1 <= lengths_104;
            end else if (8'h67 == characterIndex) begin
              lengthsOut_1 <= lengths_103;
            end else if (8'h66 == characterIndex) begin
              lengthsOut_1 <= lengths_102;
            end else if (8'h65 == characterIndex) begin
              lengthsOut_1 <= lengths_101;
            end else if (8'h64 == characterIndex) begin
              lengthsOut_1 <= lengths_100;
            end else if (8'h63 == characterIndex) begin
              lengthsOut_1 <= lengths_99;
            end else if (8'h62 == characterIndex) begin
              lengthsOut_1 <= lengths_98;
            end else if (8'h61 == characterIndex) begin
              lengthsOut_1 <= lengths_97;
            end else if (8'h60 == characterIndex) begin
              lengthsOut_1 <= lengths_96;
            end else if (8'h5f == characterIndex) begin
              lengthsOut_1 <= lengths_95;
            end else if (8'h5e == characterIndex) begin
              lengthsOut_1 <= lengths_94;
            end else if (8'h5d == characterIndex) begin
              lengthsOut_1 <= lengths_93;
            end else if (8'h5c == characterIndex) begin
              lengthsOut_1 <= lengths_92;
            end else if (8'h5b == characterIndex) begin
              lengthsOut_1 <= lengths_91;
            end else if (8'h5a == characterIndex) begin
              lengthsOut_1 <= lengths_90;
            end else if (8'h59 == characterIndex) begin
              lengthsOut_1 <= lengths_89;
            end else if (8'h58 == characterIndex) begin
              lengthsOut_1 <= lengths_88;
            end else if (8'h57 == characterIndex) begin
              lengthsOut_1 <= lengths_87;
            end else if (8'h56 == characterIndex) begin
              lengthsOut_1 <= lengths_86;
            end else if (8'h55 == characterIndex) begin
              lengthsOut_1 <= lengths_85;
            end else if (8'h54 == characterIndex) begin
              lengthsOut_1 <= lengths_84;
            end else if (8'h53 == characterIndex) begin
              lengthsOut_1 <= lengths_83;
            end else if (8'h52 == characterIndex) begin
              lengthsOut_1 <= lengths_82;
            end else if (8'h51 == characterIndex) begin
              lengthsOut_1 <= lengths_81;
            end else if (8'h50 == characterIndex) begin
              lengthsOut_1 <= lengths_80;
            end else if (8'h4f == characterIndex) begin
              lengthsOut_1 <= lengths_79;
            end else if (8'h4e == characterIndex) begin
              lengthsOut_1 <= lengths_78;
            end else if (8'h4d == characterIndex) begin
              lengthsOut_1 <= lengths_77;
            end else if (8'h4c == characterIndex) begin
              lengthsOut_1 <= lengths_76;
            end else if (8'h4b == characterIndex) begin
              lengthsOut_1 <= lengths_75;
            end else if (8'h4a == characterIndex) begin
              lengthsOut_1 <= lengths_74;
            end else if (8'h49 == characterIndex) begin
              lengthsOut_1 <= lengths_73;
            end else if (8'h48 == characterIndex) begin
              lengthsOut_1 <= lengths_72;
            end else if (8'h47 == characterIndex) begin
              lengthsOut_1 <= lengths_71;
            end else if (8'h46 == characterIndex) begin
              lengthsOut_1 <= lengths_70;
            end else if (8'h45 == characterIndex) begin
              lengthsOut_1 <= lengths_69;
            end else if (8'h44 == characterIndex) begin
              lengthsOut_1 <= lengths_68;
            end else if (8'h43 == characterIndex) begin
              lengthsOut_1 <= lengths_67;
            end else if (8'h42 == characterIndex) begin
              lengthsOut_1 <= lengths_66;
            end else if (8'h41 == characterIndex) begin
              lengthsOut_1 <= lengths_65;
            end else if (8'h40 == characterIndex) begin
              lengthsOut_1 <= lengths_64;
            end else if (8'h3f == characterIndex) begin
              lengthsOut_1 <= lengths_63;
            end else if (8'h3e == characterIndex) begin
              lengthsOut_1 <= lengths_62;
            end else if (8'h3d == characterIndex) begin
              lengthsOut_1 <= lengths_61;
            end else if (8'h3c == characterIndex) begin
              lengthsOut_1 <= lengths_60;
            end else if (8'h3b == characterIndex) begin
              lengthsOut_1 <= lengths_59;
            end else if (8'h3a == characterIndex) begin
              lengthsOut_1 <= lengths_58;
            end else if (8'h39 == characterIndex) begin
              lengthsOut_1 <= lengths_57;
            end else if (8'h38 == characterIndex) begin
              lengthsOut_1 <= lengths_56;
            end else if (8'h37 == characterIndex) begin
              lengthsOut_1 <= lengths_55;
            end else if (8'h36 == characterIndex) begin
              lengthsOut_1 <= lengths_54;
            end else if (8'h35 == characterIndex) begin
              lengthsOut_1 <= lengths_53;
            end else if (8'h34 == characterIndex) begin
              lengthsOut_1 <= lengths_52;
            end else if (8'h33 == characterIndex) begin
              lengthsOut_1 <= lengths_51;
            end else if (8'h32 == characterIndex) begin
              lengthsOut_1 <= lengths_50;
            end else if (8'h31 == characterIndex) begin
              lengthsOut_1 <= lengths_49;
            end else if (8'h30 == characterIndex) begin
              lengthsOut_1 <= lengths_48;
            end else if (8'h2f == characterIndex) begin
              lengthsOut_1 <= lengths_47;
            end else if (8'h2e == characterIndex) begin
              lengthsOut_1 <= lengths_46;
            end else if (8'h2d == characterIndex) begin
              lengthsOut_1 <= lengths_45;
            end else if (8'h2c == characterIndex) begin
              lengthsOut_1 <= lengths_44;
            end else if (8'h2b == characterIndex) begin
              lengthsOut_1 <= lengths_43;
            end else if (8'h2a == characterIndex) begin
              lengthsOut_1 <= lengths_42;
            end else if (8'h29 == characterIndex) begin
              lengthsOut_1 <= lengths_41;
            end else if (8'h28 == characterIndex) begin
              lengthsOut_1 <= lengths_40;
            end else if (8'h27 == characterIndex) begin
              lengthsOut_1 <= lengths_39;
            end else if (8'h26 == characterIndex) begin
              lengthsOut_1 <= lengths_38;
            end else if (8'h25 == characterIndex) begin
              lengthsOut_1 <= lengths_37;
            end else if (8'h24 == characterIndex) begin
              lengthsOut_1 <= lengths_36;
            end else if (8'h23 == characterIndex) begin
              lengthsOut_1 <= lengths_35;
            end else if (8'h22 == characterIndex) begin
              lengthsOut_1 <= lengths_34;
            end else if (8'h21 == characterIndex) begin
              lengthsOut_1 <= lengths_33;
            end else if (8'h20 == characterIndex) begin
              lengthsOut_1 <= lengths_32;
            end else if (8'h1f == characterIndex) begin
              lengthsOut_1 <= lengths_31;
            end else if (8'h1e == characterIndex) begin
              lengthsOut_1 <= lengths_30;
            end else if (8'h1d == characterIndex) begin
              lengthsOut_1 <= lengths_29;
            end else if (8'h1c == characterIndex) begin
              lengthsOut_1 <= lengths_28;
            end else if (8'h1b == characterIndex) begin
              lengthsOut_1 <= lengths_27;
            end else if (8'h1a == characterIndex) begin
              lengthsOut_1 <= lengths_26;
            end else if (8'h19 == characterIndex) begin
              lengthsOut_1 <= lengths_25;
            end else if (8'h18 == characterIndex) begin
              lengthsOut_1 <= lengths_24;
            end else if (8'h17 == characterIndex) begin
              lengthsOut_1 <= lengths_23;
            end else if (8'h16 == characterIndex) begin
              lengthsOut_1 <= lengths_22;
            end else if (8'h15 == characterIndex) begin
              lengthsOut_1 <= lengths_21;
            end else if (8'h14 == characterIndex) begin
              lengthsOut_1 <= lengths_20;
            end else if (8'h13 == characterIndex) begin
              lengthsOut_1 <= lengths_19;
            end else if (8'h12 == characterIndex) begin
              lengthsOut_1 <= lengths_18;
            end else if (8'h11 == characterIndex) begin
              lengthsOut_1 <= lengths_17;
            end else if (8'h10 == characterIndex) begin
              lengthsOut_1 <= lengths_16;
            end else if (8'hf == characterIndex) begin
              lengthsOut_1 <= lengths_15;
            end else if (8'he == characterIndex) begin
              lengthsOut_1 <= lengths_14;
            end else if (8'hd == characterIndex) begin
              lengthsOut_1 <= lengths_13;
            end else if (8'hc == characterIndex) begin
              lengthsOut_1 <= lengths_12;
            end else if (8'hb == characterIndex) begin
              lengthsOut_1 <= lengths_11;
            end else if (8'ha == characterIndex) begin
              lengthsOut_1 <= lengths_10;
            end else if (8'h9 == characterIndex) begin
              lengthsOut_1 <= lengths_9;
            end else if (8'h8 == characterIndex) begin
              lengthsOut_1 <= lengths_8;
            end else if (8'h7 == characterIndex) begin
              lengthsOut_1 <= lengths_7;
            end else if (8'h6 == characterIndex) begin
              lengthsOut_1 <= lengths_6;
            end else if (8'h5 == characterIndex) begin
              lengthsOut_1 <= lengths_5;
            end else if (8'h4 == characterIndex) begin
              lengthsOut_1 <= lengths_4;
            end else if (8'h3 == characterIndex) begin
              lengthsOut_1 <= lengths_3;
            end else if (8'h2 == characterIndex) begin
              lengthsOut_1 <= lengths_2;
            end else if (8'h1 == characterIndex) begin
              lengthsOut_1 <= lengths_1;
            end else begin
              lengthsOut_1 <= lengths_0;
            end
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h2 == characterIndex) begin
              lengthsOut_2 <= _T_69;
            end
          end else if (8'h2 == characterIndex) begin
            if (8'hff == characterIndex) begin
              lengthsOut_2 <= lengths_255;
            end else if (8'hfe == characterIndex) begin
              lengthsOut_2 <= lengths_254;
            end else if (8'hfd == characterIndex) begin
              lengthsOut_2 <= lengths_253;
            end else if (8'hfc == characterIndex) begin
              lengthsOut_2 <= lengths_252;
            end else if (8'hfb == characterIndex) begin
              lengthsOut_2 <= lengths_251;
            end else if (8'hfa == characterIndex) begin
              lengthsOut_2 <= lengths_250;
            end else if (8'hf9 == characterIndex) begin
              lengthsOut_2 <= lengths_249;
            end else if (8'hf8 == characterIndex) begin
              lengthsOut_2 <= lengths_248;
            end else if (8'hf7 == characterIndex) begin
              lengthsOut_2 <= lengths_247;
            end else if (8'hf6 == characterIndex) begin
              lengthsOut_2 <= lengths_246;
            end else if (8'hf5 == characterIndex) begin
              lengthsOut_2 <= lengths_245;
            end else if (8'hf4 == characterIndex) begin
              lengthsOut_2 <= lengths_244;
            end else if (8'hf3 == characterIndex) begin
              lengthsOut_2 <= lengths_243;
            end else if (8'hf2 == characterIndex) begin
              lengthsOut_2 <= lengths_242;
            end else if (8'hf1 == characterIndex) begin
              lengthsOut_2 <= lengths_241;
            end else if (8'hf0 == characterIndex) begin
              lengthsOut_2 <= lengths_240;
            end else if (8'hef == characterIndex) begin
              lengthsOut_2 <= lengths_239;
            end else if (8'hee == characterIndex) begin
              lengthsOut_2 <= lengths_238;
            end else if (8'hed == characterIndex) begin
              lengthsOut_2 <= lengths_237;
            end else if (8'hec == characterIndex) begin
              lengthsOut_2 <= lengths_236;
            end else if (8'heb == characterIndex) begin
              lengthsOut_2 <= lengths_235;
            end else if (8'hea == characterIndex) begin
              lengthsOut_2 <= lengths_234;
            end else if (8'he9 == characterIndex) begin
              lengthsOut_2 <= lengths_233;
            end else if (8'he8 == characterIndex) begin
              lengthsOut_2 <= lengths_232;
            end else if (8'he7 == characterIndex) begin
              lengthsOut_2 <= lengths_231;
            end else if (8'he6 == characterIndex) begin
              lengthsOut_2 <= lengths_230;
            end else if (8'he5 == characterIndex) begin
              lengthsOut_2 <= lengths_229;
            end else if (8'he4 == characterIndex) begin
              lengthsOut_2 <= lengths_228;
            end else if (8'he3 == characterIndex) begin
              lengthsOut_2 <= lengths_227;
            end else if (8'he2 == characterIndex) begin
              lengthsOut_2 <= lengths_226;
            end else if (8'he1 == characterIndex) begin
              lengthsOut_2 <= lengths_225;
            end else if (8'he0 == characterIndex) begin
              lengthsOut_2 <= lengths_224;
            end else if (8'hdf == characterIndex) begin
              lengthsOut_2 <= lengths_223;
            end else if (8'hde == characterIndex) begin
              lengthsOut_2 <= lengths_222;
            end else if (8'hdd == characterIndex) begin
              lengthsOut_2 <= lengths_221;
            end else if (8'hdc == characterIndex) begin
              lengthsOut_2 <= lengths_220;
            end else if (8'hdb == characterIndex) begin
              lengthsOut_2 <= lengths_219;
            end else if (8'hda == characterIndex) begin
              lengthsOut_2 <= lengths_218;
            end else if (8'hd9 == characterIndex) begin
              lengthsOut_2 <= lengths_217;
            end else if (8'hd8 == characterIndex) begin
              lengthsOut_2 <= lengths_216;
            end else if (8'hd7 == characterIndex) begin
              lengthsOut_2 <= lengths_215;
            end else if (8'hd6 == characterIndex) begin
              lengthsOut_2 <= lengths_214;
            end else if (8'hd5 == characterIndex) begin
              lengthsOut_2 <= lengths_213;
            end else if (8'hd4 == characterIndex) begin
              lengthsOut_2 <= lengths_212;
            end else if (8'hd3 == characterIndex) begin
              lengthsOut_2 <= lengths_211;
            end else if (8'hd2 == characterIndex) begin
              lengthsOut_2 <= lengths_210;
            end else if (8'hd1 == characterIndex) begin
              lengthsOut_2 <= lengths_209;
            end else if (8'hd0 == characterIndex) begin
              lengthsOut_2 <= lengths_208;
            end else if (8'hcf == characterIndex) begin
              lengthsOut_2 <= lengths_207;
            end else if (8'hce == characterIndex) begin
              lengthsOut_2 <= lengths_206;
            end else if (8'hcd == characterIndex) begin
              lengthsOut_2 <= lengths_205;
            end else if (8'hcc == characterIndex) begin
              lengthsOut_2 <= lengths_204;
            end else if (8'hcb == characterIndex) begin
              lengthsOut_2 <= lengths_203;
            end else if (8'hca == characterIndex) begin
              lengthsOut_2 <= lengths_202;
            end else if (8'hc9 == characterIndex) begin
              lengthsOut_2 <= lengths_201;
            end else if (8'hc8 == characterIndex) begin
              lengthsOut_2 <= lengths_200;
            end else if (8'hc7 == characterIndex) begin
              lengthsOut_2 <= lengths_199;
            end else if (8'hc6 == characterIndex) begin
              lengthsOut_2 <= lengths_198;
            end else if (8'hc5 == characterIndex) begin
              lengthsOut_2 <= lengths_197;
            end else if (8'hc4 == characterIndex) begin
              lengthsOut_2 <= lengths_196;
            end else if (8'hc3 == characterIndex) begin
              lengthsOut_2 <= lengths_195;
            end else if (8'hc2 == characterIndex) begin
              lengthsOut_2 <= lengths_194;
            end else if (8'hc1 == characterIndex) begin
              lengthsOut_2 <= lengths_193;
            end else if (8'hc0 == characterIndex) begin
              lengthsOut_2 <= lengths_192;
            end else if (8'hbf == characterIndex) begin
              lengthsOut_2 <= lengths_191;
            end else if (8'hbe == characterIndex) begin
              lengthsOut_2 <= lengths_190;
            end else if (8'hbd == characterIndex) begin
              lengthsOut_2 <= lengths_189;
            end else if (8'hbc == characterIndex) begin
              lengthsOut_2 <= lengths_188;
            end else if (8'hbb == characterIndex) begin
              lengthsOut_2 <= lengths_187;
            end else if (8'hba == characterIndex) begin
              lengthsOut_2 <= lengths_186;
            end else if (8'hb9 == characterIndex) begin
              lengthsOut_2 <= lengths_185;
            end else if (8'hb8 == characterIndex) begin
              lengthsOut_2 <= lengths_184;
            end else if (8'hb7 == characterIndex) begin
              lengthsOut_2 <= lengths_183;
            end else if (8'hb6 == characterIndex) begin
              lengthsOut_2 <= lengths_182;
            end else if (8'hb5 == characterIndex) begin
              lengthsOut_2 <= lengths_181;
            end else if (8'hb4 == characterIndex) begin
              lengthsOut_2 <= lengths_180;
            end else if (8'hb3 == characterIndex) begin
              lengthsOut_2 <= lengths_179;
            end else if (8'hb2 == characterIndex) begin
              lengthsOut_2 <= lengths_178;
            end else if (8'hb1 == characterIndex) begin
              lengthsOut_2 <= lengths_177;
            end else if (8'hb0 == characterIndex) begin
              lengthsOut_2 <= lengths_176;
            end else if (8'haf == characterIndex) begin
              lengthsOut_2 <= lengths_175;
            end else if (8'hae == characterIndex) begin
              lengthsOut_2 <= lengths_174;
            end else if (8'had == characterIndex) begin
              lengthsOut_2 <= lengths_173;
            end else if (8'hac == characterIndex) begin
              lengthsOut_2 <= lengths_172;
            end else if (8'hab == characterIndex) begin
              lengthsOut_2 <= lengths_171;
            end else if (8'haa == characterIndex) begin
              lengthsOut_2 <= lengths_170;
            end else if (8'ha9 == characterIndex) begin
              lengthsOut_2 <= lengths_169;
            end else if (8'ha8 == characterIndex) begin
              lengthsOut_2 <= lengths_168;
            end else if (8'ha7 == characterIndex) begin
              lengthsOut_2 <= lengths_167;
            end else if (8'ha6 == characterIndex) begin
              lengthsOut_2 <= lengths_166;
            end else if (8'ha5 == characterIndex) begin
              lengthsOut_2 <= lengths_165;
            end else if (8'ha4 == characterIndex) begin
              lengthsOut_2 <= lengths_164;
            end else if (8'ha3 == characterIndex) begin
              lengthsOut_2 <= lengths_163;
            end else if (8'ha2 == characterIndex) begin
              lengthsOut_2 <= lengths_162;
            end else if (8'ha1 == characterIndex) begin
              lengthsOut_2 <= lengths_161;
            end else if (8'ha0 == characterIndex) begin
              lengthsOut_2 <= lengths_160;
            end else if (8'h9f == characterIndex) begin
              lengthsOut_2 <= lengths_159;
            end else if (8'h9e == characterIndex) begin
              lengthsOut_2 <= lengths_158;
            end else if (8'h9d == characterIndex) begin
              lengthsOut_2 <= lengths_157;
            end else if (8'h9c == characterIndex) begin
              lengthsOut_2 <= lengths_156;
            end else if (8'h9b == characterIndex) begin
              lengthsOut_2 <= lengths_155;
            end else if (8'h9a == characterIndex) begin
              lengthsOut_2 <= lengths_154;
            end else if (8'h99 == characterIndex) begin
              lengthsOut_2 <= lengths_153;
            end else if (8'h98 == characterIndex) begin
              lengthsOut_2 <= lengths_152;
            end else if (8'h97 == characterIndex) begin
              lengthsOut_2 <= lengths_151;
            end else if (8'h96 == characterIndex) begin
              lengthsOut_2 <= lengths_150;
            end else if (8'h95 == characterIndex) begin
              lengthsOut_2 <= lengths_149;
            end else if (8'h94 == characterIndex) begin
              lengthsOut_2 <= lengths_148;
            end else if (8'h93 == characterIndex) begin
              lengthsOut_2 <= lengths_147;
            end else if (8'h92 == characterIndex) begin
              lengthsOut_2 <= lengths_146;
            end else if (8'h91 == characterIndex) begin
              lengthsOut_2 <= lengths_145;
            end else if (8'h90 == characterIndex) begin
              lengthsOut_2 <= lengths_144;
            end else if (8'h8f == characterIndex) begin
              lengthsOut_2 <= lengths_143;
            end else if (8'h8e == characterIndex) begin
              lengthsOut_2 <= lengths_142;
            end else if (8'h8d == characterIndex) begin
              lengthsOut_2 <= lengths_141;
            end else if (8'h8c == characterIndex) begin
              lengthsOut_2 <= lengths_140;
            end else if (8'h8b == characterIndex) begin
              lengthsOut_2 <= lengths_139;
            end else if (8'h8a == characterIndex) begin
              lengthsOut_2 <= lengths_138;
            end else if (8'h89 == characterIndex) begin
              lengthsOut_2 <= lengths_137;
            end else if (8'h88 == characterIndex) begin
              lengthsOut_2 <= lengths_136;
            end else if (8'h87 == characterIndex) begin
              lengthsOut_2 <= lengths_135;
            end else if (8'h86 == characterIndex) begin
              lengthsOut_2 <= lengths_134;
            end else if (8'h85 == characterIndex) begin
              lengthsOut_2 <= lengths_133;
            end else if (8'h84 == characterIndex) begin
              lengthsOut_2 <= lengths_132;
            end else if (8'h83 == characterIndex) begin
              lengthsOut_2 <= lengths_131;
            end else if (8'h82 == characterIndex) begin
              lengthsOut_2 <= lengths_130;
            end else if (8'h81 == characterIndex) begin
              lengthsOut_2 <= lengths_129;
            end else if (8'h80 == characterIndex) begin
              lengthsOut_2 <= lengths_128;
            end else if (8'h7f == characterIndex) begin
              lengthsOut_2 <= lengths_127;
            end else if (8'h7e == characterIndex) begin
              lengthsOut_2 <= lengths_126;
            end else if (8'h7d == characterIndex) begin
              lengthsOut_2 <= lengths_125;
            end else if (8'h7c == characterIndex) begin
              lengthsOut_2 <= lengths_124;
            end else if (8'h7b == characterIndex) begin
              lengthsOut_2 <= lengths_123;
            end else if (8'h7a == characterIndex) begin
              lengthsOut_2 <= lengths_122;
            end else if (8'h79 == characterIndex) begin
              lengthsOut_2 <= lengths_121;
            end else if (8'h78 == characterIndex) begin
              lengthsOut_2 <= lengths_120;
            end else if (8'h77 == characterIndex) begin
              lengthsOut_2 <= lengths_119;
            end else if (8'h76 == characterIndex) begin
              lengthsOut_2 <= lengths_118;
            end else if (8'h75 == characterIndex) begin
              lengthsOut_2 <= lengths_117;
            end else if (8'h74 == characterIndex) begin
              lengthsOut_2 <= lengths_116;
            end else if (8'h73 == characterIndex) begin
              lengthsOut_2 <= lengths_115;
            end else if (8'h72 == characterIndex) begin
              lengthsOut_2 <= lengths_114;
            end else if (8'h71 == characterIndex) begin
              lengthsOut_2 <= lengths_113;
            end else if (8'h70 == characterIndex) begin
              lengthsOut_2 <= lengths_112;
            end else if (8'h6f == characterIndex) begin
              lengthsOut_2 <= lengths_111;
            end else if (8'h6e == characterIndex) begin
              lengthsOut_2 <= lengths_110;
            end else if (8'h6d == characterIndex) begin
              lengthsOut_2 <= lengths_109;
            end else if (8'h6c == characterIndex) begin
              lengthsOut_2 <= lengths_108;
            end else if (8'h6b == characterIndex) begin
              lengthsOut_2 <= lengths_107;
            end else if (8'h6a == characterIndex) begin
              lengthsOut_2 <= lengths_106;
            end else if (8'h69 == characterIndex) begin
              lengthsOut_2 <= lengths_105;
            end else if (8'h68 == characterIndex) begin
              lengthsOut_2 <= lengths_104;
            end else if (8'h67 == characterIndex) begin
              lengthsOut_2 <= lengths_103;
            end else if (8'h66 == characterIndex) begin
              lengthsOut_2 <= lengths_102;
            end else if (8'h65 == characterIndex) begin
              lengthsOut_2 <= lengths_101;
            end else if (8'h64 == characterIndex) begin
              lengthsOut_2 <= lengths_100;
            end else if (8'h63 == characterIndex) begin
              lengthsOut_2 <= lengths_99;
            end else if (8'h62 == characterIndex) begin
              lengthsOut_2 <= lengths_98;
            end else if (8'h61 == characterIndex) begin
              lengthsOut_2 <= lengths_97;
            end else if (8'h60 == characterIndex) begin
              lengthsOut_2 <= lengths_96;
            end else if (8'h5f == characterIndex) begin
              lengthsOut_2 <= lengths_95;
            end else if (8'h5e == characterIndex) begin
              lengthsOut_2 <= lengths_94;
            end else if (8'h5d == characterIndex) begin
              lengthsOut_2 <= lengths_93;
            end else if (8'h5c == characterIndex) begin
              lengthsOut_2 <= lengths_92;
            end else if (8'h5b == characterIndex) begin
              lengthsOut_2 <= lengths_91;
            end else if (8'h5a == characterIndex) begin
              lengthsOut_2 <= lengths_90;
            end else if (8'h59 == characterIndex) begin
              lengthsOut_2 <= lengths_89;
            end else if (8'h58 == characterIndex) begin
              lengthsOut_2 <= lengths_88;
            end else if (8'h57 == characterIndex) begin
              lengthsOut_2 <= lengths_87;
            end else if (8'h56 == characterIndex) begin
              lengthsOut_2 <= lengths_86;
            end else if (8'h55 == characterIndex) begin
              lengthsOut_2 <= lengths_85;
            end else if (8'h54 == characterIndex) begin
              lengthsOut_2 <= lengths_84;
            end else if (8'h53 == characterIndex) begin
              lengthsOut_2 <= lengths_83;
            end else if (8'h52 == characterIndex) begin
              lengthsOut_2 <= lengths_82;
            end else if (8'h51 == characterIndex) begin
              lengthsOut_2 <= lengths_81;
            end else if (8'h50 == characterIndex) begin
              lengthsOut_2 <= lengths_80;
            end else if (8'h4f == characterIndex) begin
              lengthsOut_2 <= lengths_79;
            end else if (8'h4e == characterIndex) begin
              lengthsOut_2 <= lengths_78;
            end else if (8'h4d == characterIndex) begin
              lengthsOut_2 <= lengths_77;
            end else if (8'h4c == characterIndex) begin
              lengthsOut_2 <= lengths_76;
            end else if (8'h4b == characterIndex) begin
              lengthsOut_2 <= lengths_75;
            end else if (8'h4a == characterIndex) begin
              lengthsOut_2 <= lengths_74;
            end else if (8'h49 == characterIndex) begin
              lengthsOut_2 <= lengths_73;
            end else if (8'h48 == characterIndex) begin
              lengthsOut_2 <= lengths_72;
            end else if (8'h47 == characterIndex) begin
              lengthsOut_2 <= lengths_71;
            end else if (8'h46 == characterIndex) begin
              lengthsOut_2 <= lengths_70;
            end else if (8'h45 == characterIndex) begin
              lengthsOut_2 <= lengths_69;
            end else if (8'h44 == characterIndex) begin
              lengthsOut_2 <= lengths_68;
            end else if (8'h43 == characterIndex) begin
              lengthsOut_2 <= lengths_67;
            end else if (8'h42 == characterIndex) begin
              lengthsOut_2 <= lengths_66;
            end else if (8'h41 == characterIndex) begin
              lengthsOut_2 <= lengths_65;
            end else if (8'h40 == characterIndex) begin
              lengthsOut_2 <= lengths_64;
            end else if (8'h3f == characterIndex) begin
              lengthsOut_2 <= lengths_63;
            end else if (8'h3e == characterIndex) begin
              lengthsOut_2 <= lengths_62;
            end else if (8'h3d == characterIndex) begin
              lengthsOut_2 <= lengths_61;
            end else if (8'h3c == characterIndex) begin
              lengthsOut_2 <= lengths_60;
            end else if (8'h3b == characterIndex) begin
              lengthsOut_2 <= lengths_59;
            end else if (8'h3a == characterIndex) begin
              lengthsOut_2 <= lengths_58;
            end else if (8'h39 == characterIndex) begin
              lengthsOut_2 <= lengths_57;
            end else if (8'h38 == characterIndex) begin
              lengthsOut_2 <= lengths_56;
            end else if (8'h37 == characterIndex) begin
              lengthsOut_2 <= lengths_55;
            end else if (8'h36 == characterIndex) begin
              lengthsOut_2 <= lengths_54;
            end else if (8'h35 == characterIndex) begin
              lengthsOut_2 <= lengths_53;
            end else if (8'h34 == characterIndex) begin
              lengthsOut_2 <= lengths_52;
            end else if (8'h33 == characterIndex) begin
              lengthsOut_2 <= lengths_51;
            end else if (8'h32 == characterIndex) begin
              lengthsOut_2 <= lengths_50;
            end else if (8'h31 == characterIndex) begin
              lengthsOut_2 <= lengths_49;
            end else if (8'h30 == characterIndex) begin
              lengthsOut_2 <= lengths_48;
            end else if (8'h2f == characterIndex) begin
              lengthsOut_2 <= lengths_47;
            end else if (8'h2e == characterIndex) begin
              lengthsOut_2 <= lengths_46;
            end else if (8'h2d == characterIndex) begin
              lengthsOut_2 <= lengths_45;
            end else if (8'h2c == characterIndex) begin
              lengthsOut_2 <= lengths_44;
            end else if (8'h2b == characterIndex) begin
              lengthsOut_2 <= lengths_43;
            end else if (8'h2a == characterIndex) begin
              lengthsOut_2 <= lengths_42;
            end else if (8'h29 == characterIndex) begin
              lengthsOut_2 <= lengths_41;
            end else if (8'h28 == characterIndex) begin
              lengthsOut_2 <= lengths_40;
            end else if (8'h27 == characterIndex) begin
              lengthsOut_2 <= lengths_39;
            end else if (8'h26 == characterIndex) begin
              lengthsOut_2 <= lengths_38;
            end else if (8'h25 == characterIndex) begin
              lengthsOut_2 <= lengths_37;
            end else if (8'h24 == characterIndex) begin
              lengthsOut_2 <= lengths_36;
            end else if (8'h23 == characterIndex) begin
              lengthsOut_2 <= lengths_35;
            end else if (8'h22 == characterIndex) begin
              lengthsOut_2 <= lengths_34;
            end else if (8'h21 == characterIndex) begin
              lengthsOut_2 <= lengths_33;
            end else if (8'h20 == characterIndex) begin
              lengthsOut_2 <= lengths_32;
            end else if (8'h1f == characterIndex) begin
              lengthsOut_2 <= lengths_31;
            end else if (8'h1e == characterIndex) begin
              lengthsOut_2 <= lengths_30;
            end else if (8'h1d == characterIndex) begin
              lengthsOut_2 <= lengths_29;
            end else if (8'h1c == characterIndex) begin
              lengthsOut_2 <= lengths_28;
            end else if (8'h1b == characterIndex) begin
              lengthsOut_2 <= lengths_27;
            end else if (8'h1a == characterIndex) begin
              lengthsOut_2 <= lengths_26;
            end else if (8'h19 == characterIndex) begin
              lengthsOut_2 <= lengths_25;
            end else if (8'h18 == characterIndex) begin
              lengthsOut_2 <= lengths_24;
            end else if (8'h17 == characterIndex) begin
              lengthsOut_2 <= lengths_23;
            end else if (8'h16 == characterIndex) begin
              lengthsOut_2 <= lengths_22;
            end else if (8'h15 == characterIndex) begin
              lengthsOut_2 <= lengths_21;
            end else if (8'h14 == characterIndex) begin
              lengthsOut_2 <= lengths_20;
            end else if (8'h13 == characterIndex) begin
              lengthsOut_2 <= lengths_19;
            end else if (8'h12 == characterIndex) begin
              lengthsOut_2 <= lengths_18;
            end else if (8'h11 == characterIndex) begin
              lengthsOut_2 <= lengths_17;
            end else if (8'h10 == characterIndex) begin
              lengthsOut_2 <= lengths_16;
            end else if (8'hf == characterIndex) begin
              lengthsOut_2 <= lengths_15;
            end else if (8'he == characterIndex) begin
              lengthsOut_2 <= lengths_14;
            end else if (8'hd == characterIndex) begin
              lengthsOut_2 <= lengths_13;
            end else if (8'hc == characterIndex) begin
              lengthsOut_2 <= lengths_12;
            end else if (8'hb == characterIndex) begin
              lengthsOut_2 <= lengths_11;
            end else if (8'ha == characterIndex) begin
              lengthsOut_2 <= lengths_10;
            end else if (8'h9 == characterIndex) begin
              lengthsOut_2 <= lengths_9;
            end else if (8'h8 == characterIndex) begin
              lengthsOut_2 <= lengths_8;
            end else if (8'h7 == characterIndex) begin
              lengthsOut_2 <= lengths_7;
            end else if (8'h6 == characterIndex) begin
              lengthsOut_2 <= lengths_6;
            end else if (8'h5 == characterIndex) begin
              lengthsOut_2 <= lengths_5;
            end else if (8'h4 == characterIndex) begin
              lengthsOut_2 <= lengths_4;
            end else if (8'h3 == characterIndex) begin
              lengthsOut_2 <= lengths_3;
            end else if (8'h2 == characterIndex) begin
              lengthsOut_2 <= lengths_2;
            end else if (8'h1 == characterIndex) begin
              lengthsOut_2 <= lengths_1;
            end else begin
              lengthsOut_2 <= lengths_0;
            end
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h3 == characterIndex) begin
              lengthsOut_3 <= _T_69;
            end
          end else if (8'h3 == characterIndex) begin
            if (8'hff == characterIndex) begin
              lengthsOut_3 <= lengths_255;
            end else if (8'hfe == characterIndex) begin
              lengthsOut_3 <= lengths_254;
            end else if (8'hfd == characterIndex) begin
              lengthsOut_3 <= lengths_253;
            end else if (8'hfc == characterIndex) begin
              lengthsOut_3 <= lengths_252;
            end else if (8'hfb == characterIndex) begin
              lengthsOut_3 <= lengths_251;
            end else if (8'hfa == characterIndex) begin
              lengthsOut_3 <= lengths_250;
            end else if (8'hf9 == characterIndex) begin
              lengthsOut_3 <= lengths_249;
            end else if (8'hf8 == characterIndex) begin
              lengthsOut_3 <= lengths_248;
            end else if (8'hf7 == characterIndex) begin
              lengthsOut_3 <= lengths_247;
            end else if (8'hf6 == characterIndex) begin
              lengthsOut_3 <= lengths_246;
            end else if (8'hf5 == characterIndex) begin
              lengthsOut_3 <= lengths_245;
            end else if (8'hf4 == characterIndex) begin
              lengthsOut_3 <= lengths_244;
            end else if (8'hf3 == characterIndex) begin
              lengthsOut_3 <= lengths_243;
            end else if (8'hf2 == characterIndex) begin
              lengthsOut_3 <= lengths_242;
            end else if (8'hf1 == characterIndex) begin
              lengthsOut_3 <= lengths_241;
            end else if (8'hf0 == characterIndex) begin
              lengthsOut_3 <= lengths_240;
            end else if (8'hef == characterIndex) begin
              lengthsOut_3 <= lengths_239;
            end else if (8'hee == characterIndex) begin
              lengthsOut_3 <= lengths_238;
            end else if (8'hed == characterIndex) begin
              lengthsOut_3 <= lengths_237;
            end else if (8'hec == characterIndex) begin
              lengthsOut_3 <= lengths_236;
            end else if (8'heb == characterIndex) begin
              lengthsOut_3 <= lengths_235;
            end else if (8'hea == characterIndex) begin
              lengthsOut_3 <= lengths_234;
            end else if (8'he9 == characterIndex) begin
              lengthsOut_3 <= lengths_233;
            end else if (8'he8 == characterIndex) begin
              lengthsOut_3 <= lengths_232;
            end else if (8'he7 == characterIndex) begin
              lengthsOut_3 <= lengths_231;
            end else if (8'he6 == characterIndex) begin
              lengthsOut_3 <= lengths_230;
            end else if (8'he5 == characterIndex) begin
              lengthsOut_3 <= lengths_229;
            end else if (8'he4 == characterIndex) begin
              lengthsOut_3 <= lengths_228;
            end else if (8'he3 == characterIndex) begin
              lengthsOut_3 <= lengths_227;
            end else if (8'he2 == characterIndex) begin
              lengthsOut_3 <= lengths_226;
            end else if (8'he1 == characterIndex) begin
              lengthsOut_3 <= lengths_225;
            end else if (8'he0 == characterIndex) begin
              lengthsOut_3 <= lengths_224;
            end else if (8'hdf == characterIndex) begin
              lengthsOut_3 <= lengths_223;
            end else if (8'hde == characterIndex) begin
              lengthsOut_3 <= lengths_222;
            end else if (8'hdd == characterIndex) begin
              lengthsOut_3 <= lengths_221;
            end else if (8'hdc == characterIndex) begin
              lengthsOut_3 <= lengths_220;
            end else if (8'hdb == characterIndex) begin
              lengthsOut_3 <= lengths_219;
            end else if (8'hda == characterIndex) begin
              lengthsOut_3 <= lengths_218;
            end else if (8'hd9 == characterIndex) begin
              lengthsOut_3 <= lengths_217;
            end else if (8'hd8 == characterIndex) begin
              lengthsOut_3 <= lengths_216;
            end else if (8'hd7 == characterIndex) begin
              lengthsOut_3 <= lengths_215;
            end else if (8'hd6 == characterIndex) begin
              lengthsOut_3 <= lengths_214;
            end else if (8'hd5 == characterIndex) begin
              lengthsOut_3 <= lengths_213;
            end else if (8'hd4 == characterIndex) begin
              lengthsOut_3 <= lengths_212;
            end else if (8'hd3 == characterIndex) begin
              lengthsOut_3 <= lengths_211;
            end else if (8'hd2 == characterIndex) begin
              lengthsOut_3 <= lengths_210;
            end else if (8'hd1 == characterIndex) begin
              lengthsOut_3 <= lengths_209;
            end else if (8'hd0 == characterIndex) begin
              lengthsOut_3 <= lengths_208;
            end else if (8'hcf == characterIndex) begin
              lengthsOut_3 <= lengths_207;
            end else if (8'hce == characterIndex) begin
              lengthsOut_3 <= lengths_206;
            end else if (8'hcd == characterIndex) begin
              lengthsOut_3 <= lengths_205;
            end else if (8'hcc == characterIndex) begin
              lengthsOut_3 <= lengths_204;
            end else if (8'hcb == characterIndex) begin
              lengthsOut_3 <= lengths_203;
            end else if (8'hca == characterIndex) begin
              lengthsOut_3 <= lengths_202;
            end else if (8'hc9 == characterIndex) begin
              lengthsOut_3 <= lengths_201;
            end else if (8'hc8 == characterIndex) begin
              lengthsOut_3 <= lengths_200;
            end else if (8'hc7 == characterIndex) begin
              lengthsOut_3 <= lengths_199;
            end else if (8'hc6 == characterIndex) begin
              lengthsOut_3 <= lengths_198;
            end else if (8'hc5 == characterIndex) begin
              lengthsOut_3 <= lengths_197;
            end else if (8'hc4 == characterIndex) begin
              lengthsOut_3 <= lengths_196;
            end else if (8'hc3 == characterIndex) begin
              lengthsOut_3 <= lengths_195;
            end else if (8'hc2 == characterIndex) begin
              lengthsOut_3 <= lengths_194;
            end else if (8'hc1 == characterIndex) begin
              lengthsOut_3 <= lengths_193;
            end else if (8'hc0 == characterIndex) begin
              lengthsOut_3 <= lengths_192;
            end else if (8'hbf == characterIndex) begin
              lengthsOut_3 <= lengths_191;
            end else if (8'hbe == characterIndex) begin
              lengthsOut_3 <= lengths_190;
            end else if (8'hbd == characterIndex) begin
              lengthsOut_3 <= lengths_189;
            end else if (8'hbc == characterIndex) begin
              lengthsOut_3 <= lengths_188;
            end else if (8'hbb == characterIndex) begin
              lengthsOut_3 <= lengths_187;
            end else if (8'hba == characterIndex) begin
              lengthsOut_3 <= lengths_186;
            end else if (8'hb9 == characterIndex) begin
              lengthsOut_3 <= lengths_185;
            end else if (8'hb8 == characterIndex) begin
              lengthsOut_3 <= lengths_184;
            end else if (8'hb7 == characterIndex) begin
              lengthsOut_3 <= lengths_183;
            end else if (8'hb6 == characterIndex) begin
              lengthsOut_3 <= lengths_182;
            end else if (8'hb5 == characterIndex) begin
              lengthsOut_3 <= lengths_181;
            end else if (8'hb4 == characterIndex) begin
              lengthsOut_3 <= lengths_180;
            end else if (8'hb3 == characterIndex) begin
              lengthsOut_3 <= lengths_179;
            end else if (8'hb2 == characterIndex) begin
              lengthsOut_3 <= lengths_178;
            end else if (8'hb1 == characterIndex) begin
              lengthsOut_3 <= lengths_177;
            end else if (8'hb0 == characterIndex) begin
              lengthsOut_3 <= lengths_176;
            end else if (8'haf == characterIndex) begin
              lengthsOut_3 <= lengths_175;
            end else if (8'hae == characterIndex) begin
              lengthsOut_3 <= lengths_174;
            end else if (8'had == characterIndex) begin
              lengthsOut_3 <= lengths_173;
            end else if (8'hac == characterIndex) begin
              lengthsOut_3 <= lengths_172;
            end else if (8'hab == characterIndex) begin
              lengthsOut_3 <= lengths_171;
            end else if (8'haa == characterIndex) begin
              lengthsOut_3 <= lengths_170;
            end else if (8'ha9 == characterIndex) begin
              lengthsOut_3 <= lengths_169;
            end else if (8'ha8 == characterIndex) begin
              lengthsOut_3 <= lengths_168;
            end else if (8'ha7 == characterIndex) begin
              lengthsOut_3 <= lengths_167;
            end else if (8'ha6 == characterIndex) begin
              lengthsOut_3 <= lengths_166;
            end else if (8'ha5 == characterIndex) begin
              lengthsOut_3 <= lengths_165;
            end else if (8'ha4 == characterIndex) begin
              lengthsOut_3 <= lengths_164;
            end else if (8'ha3 == characterIndex) begin
              lengthsOut_3 <= lengths_163;
            end else if (8'ha2 == characterIndex) begin
              lengthsOut_3 <= lengths_162;
            end else if (8'ha1 == characterIndex) begin
              lengthsOut_3 <= lengths_161;
            end else if (8'ha0 == characterIndex) begin
              lengthsOut_3 <= lengths_160;
            end else if (8'h9f == characterIndex) begin
              lengthsOut_3 <= lengths_159;
            end else if (8'h9e == characterIndex) begin
              lengthsOut_3 <= lengths_158;
            end else if (8'h9d == characterIndex) begin
              lengthsOut_3 <= lengths_157;
            end else if (8'h9c == characterIndex) begin
              lengthsOut_3 <= lengths_156;
            end else if (8'h9b == characterIndex) begin
              lengthsOut_3 <= lengths_155;
            end else if (8'h9a == characterIndex) begin
              lengthsOut_3 <= lengths_154;
            end else if (8'h99 == characterIndex) begin
              lengthsOut_3 <= lengths_153;
            end else if (8'h98 == characterIndex) begin
              lengthsOut_3 <= lengths_152;
            end else if (8'h97 == characterIndex) begin
              lengthsOut_3 <= lengths_151;
            end else if (8'h96 == characterIndex) begin
              lengthsOut_3 <= lengths_150;
            end else if (8'h95 == characterIndex) begin
              lengthsOut_3 <= lengths_149;
            end else if (8'h94 == characterIndex) begin
              lengthsOut_3 <= lengths_148;
            end else if (8'h93 == characterIndex) begin
              lengthsOut_3 <= lengths_147;
            end else if (8'h92 == characterIndex) begin
              lengthsOut_3 <= lengths_146;
            end else if (8'h91 == characterIndex) begin
              lengthsOut_3 <= lengths_145;
            end else if (8'h90 == characterIndex) begin
              lengthsOut_3 <= lengths_144;
            end else if (8'h8f == characterIndex) begin
              lengthsOut_3 <= lengths_143;
            end else if (8'h8e == characterIndex) begin
              lengthsOut_3 <= lengths_142;
            end else if (8'h8d == characterIndex) begin
              lengthsOut_3 <= lengths_141;
            end else if (8'h8c == characterIndex) begin
              lengthsOut_3 <= lengths_140;
            end else if (8'h8b == characterIndex) begin
              lengthsOut_3 <= lengths_139;
            end else if (8'h8a == characterIndex) begin
              lengthsOut_3 <= lengths_138;
            end else if (8'h89 == characterIndex) begin
              lengthsOut_3 <= lengths_137;
            end else if (8'h88 == characterIndex) begin
              lengthsOut_3 <= lengths_136;
            end else if (8'h87 == characterIndex) begin
              lengthsOut_3 <= lengths_135;
            end else if (8'h86 == characterIndex) begin
              lengthsOut_3 <= lengths_134;
            end else if (8'h85 == characterIndex) begin
              lengthsOut_3 <= lengths_133;
            end else if (8'h84 == characterIndex) begin
              lengthsOut_3 <= lengths_132;
            end else if (8'h83 == characterIndex) begin
              lengthsOut_3 <= lengths_131;
            end else if (8'h82 == characterIndex) begin
              lengthsOut_3 <= lengths_130;
            end else if (8'h81 == characterIndex) begin
              lengthsOut_3 <= lengths_129;
            end else if (8'h80 == characterIndex) begin
              lengthsOut_3 <= lengths_128;
            end else if (8'h7f == characterIndex) begin
              lengthsOut_3 <= lengths_127;
            end else if (8'h7e == characterIndex) begin
              lengthsOut_3 <= lengths_126;
            end else if (8'h7d == characterIndex) begin
              lengthsOut_3 <= lengths_125;
            end else if (8'h7c == characterIndex) begin
              lengthsOut_3 <= lengths_124;
            end else if (8'h7b == characterIndex) begin
              lengthsOut_3 <= lengths_123;
            end else if (8'h7a == characterIndex) begin
              lengthsOut_3 <= lengths_122;
            end else if (8'h79 == characterIndex) begin
              lengthsOut_3 <= lengths_121;
            end else if (8'h78 == characterIndex) begin
              lengthsOut_3 <= lengths_120;
            end else if (8'h77 == characterIndex) begin
              lengthsOut_3 <= lengths_119;
            end else if (8'h76 == characterIndex) begin
              lengthsOut_3 <= lengths_118;
            end else if (8'h75 == characterIndex) begin
              lengthsOut_3 <= lengths_117;
            end else if (8'h74 == characterIndex) begin
              lengthsOut_3 <= lengths_116;
            end else if (8'h73 == characterIndex) begin
              lengthsOut_3 <= lengths_115;
            end else if (8'h72 == characterIndex) begin
              lengthsOut_3 <= lengths_114;
            end else if (8'h71 == characterIndex) begin
              lengthsOut_3 <= lengths_113;
            end else if (8'h70 == characterIndex) begin
              lengthsOut_3 <= lengths_112;
            end else if (8'h6f == characterIndex) begin
              lengthsOut_3 <= lengths_111;
            end else if (8'h6e == characterIndex) begin
              lengthsOut_3 <= lengths_110;
            end else if (8'h6d == characterIndex) begin
              lengthsOut_3 <= lengths_109;
            end else if (8'h6c == characterIndex) begin
              lengthsOut_3 <= lengths_108;
            end else if (8'h6b == characterIndex) begin
              lengthsOut_3 <= lengths_107;
            end else if (8'h6a == characterIndex) begin
              lengthsOut_3 <= lengths_106;
            end else if (8'h69 == characterIndex) begin
              lengthsOut_3 <= lengths_105;
            end else if (8'h68 == characterIndex) begin
              lengthsOut_3 <= lengths_104;
            end else if (8'h67 == characterIndex) begin
              lengthsOut_3 <= lengths_103;
            end else if (8'h66 == characterIndex) begin
              lengthsOut_3 <= lengths_102;
            end else if (8'h65 == characterIndex) begin
              lengthsOut_3 <= lengths_101;
            end else if (8'h64 == characterIndex) begin
              lengthsOut_3 <= lengths_100;
            end else if (8'h63 == characterIndex) begin
              lengthsOut_3 <= lengths_99;
            end else if (8'h62 == characterIndex) begin
              lengthsOut_3 <= lengths_98;
            end else if (8'h61 == characterIndex) begin
              lengthsOut_3 <= lengths_97;
            end else if (8'h60 == characterIndex) begin
              lengthsOut_3 <= lengths_96;
            end else if (8'h5f == characterIndex) begin
              lengthsOut_3 <= lengths_95;
            end else if (8'h5e == characterIndex) begin
              lengthsOut_3 <= lengths_94;
            end else if (8'h5d == characterIndex) begin
              lengthsOut_3 <= lengths_93;
            end else if (8'h5c == characterIndex) begin
              lengthsOut_3 <= lengths_92;
            end else if (8'h5b == characterIndex) begin
              lengthsOut_3 <= lengths_91;
            end else if (8'h5a == characterIndex) begin
              lengthsOut_3 <= lengths_90;
            end else if (8'h59 == characterIndex) begin
              lengthsOut_3 <= lengths_89;
            end else if (8'h58 == characterIndex) begin
              lengthsOut_3 <= lengths_88;
            end else if (8'h57 == characterIndex) begin
              lengthsOut_3 <= lengths_87;
            end else if (8'h56 == characterIndex) begin
              lengthsOut_3 <= lengths_86;
            end else if (8'h55 == characterIndex) begin
              lengthsOut_3 <= lengths_85;
            end else if (8'h54 == characterIndex) begin
              lengthsOut_3 <= lengths_84;
            end else if (8'h53 == characterIndex) begin
              lengthsOut_3 <= lengths_83;
            end else if (8'h52 == characterIndex) begin
              lengthsOut_3 <= lengths_82;
            end else if (8'h51 == characterIndex) begin
              lengthsOut_3 <= lengths_81;
            end else if (8'h50 == characterIndex) begin
              lengthsOut_3 <= lengths_80;
            end else if (8'h4f == characterIndex) begin
              lengthsOut_3 <= lengths_79;
            end else if (8'h4e == characterIndex) begin
              lengthsOut_3 <= lengths_78;
            end else if (8'h4d == characterIndex) begin
              lengthsOut_3 <= lengths_77;
            end else if (8'h4c == characterIndex) begin
              lengthsOut_3 <= lengths_76;
            end else if (8'h4b == characterIndex) begin
              lengthsOut_3 <= lengths_75;
            end else if (8'h4a == characterIndex) begin
              lengthsOut_3 <= lengths_74;
            end else if (8'h49 == characterIndex) begin
              lengthsOut_3 <= lengths_73;
            end else if (8'h48 == characterIndex) begin
              lengthsOut_3 <= lengths_72;
            end else if (8'h47 == characterIndex) begin
              lengthsOut_3 <= lengths_71;
            end else if (8'h46 == characterIndex) begin
              lengthsOut_3 <= lengths_70;
            end else if (8'h45 == characterIndex) begin
              lengthsOut_3 <= lengths_69;
            end else if (8'h44 == characterIndex) begin
              lengthsOut_3 <= lengths_68;
            end else if (8'h43 == characterIndex) begin
              lengthsOut_3 <= lengths_67;
            end else if (8'h42 == characterIndex) begin
              lengthsOut_3 <= lengths_66;
            end else if (8'h41 == characterIndex) begin
              lengthsOut_3 <= lengths_65;
            end else if (8'h40 == characterIndex) begin
              lengthsOut_3 <= lengths_64;
            end else if (8'h3f == characterIndex) begin
              lengthsOut_3 <= lengths_63;
            end else if (8'h3e == characterIndex) begin
              lengthsOut_3 <= lengths_62;
            end else if (8'h3d == characterIndex) begin
              lengthsOut_3 <= lengths_61;
            end else if (8'h3c == characterIndex) begin
              lengthsOut_3 <= lengths_60;
            end else if (8'h3b == characterIndex) begin
              lengthsOut_3 <= lengths_59;
            end else if (8'h3a == characterIndex) begin
              lengthsOut_3 <= lengths_58;
            end else if (8'h39 == characterIndex) begin
              lengthsOut_3 <= lengths_57;
            end else if (8'h38 == characterIndex) begin
              lengthsOut_3 <= lengths_56;
            end else if (8'h37 == characterIndex) begin
              lengthsOut_3 <= lengths_55;
            end else if (8'h36 == characterIndex) begin
              lengthsOut_3 <= lengths_54;
            end else if (8'h35 == characterIndex) begin
              lengthsOut_3 <= lengths_53;
            end else if (8'h34 == characterIndex) begin
              lengthsOut_3 <= lengths_52;
            end else if (8'h33 == characterIndex) begin
              lengthsOut_3 <= lengths_51;
            end else if (8'h32 == characterIndex) begin
              lengthsOut_3 <= lengths_50;
            end else if (8'h31 == characterIndex) begin
              lengthsOut_3 <= lengths_49;
            end else if (8'h30 == characterIndex) begin
              lengthsOut_3 <= lengths_48;
            end else if (8'h2f == characterIndex) begin
              lengthsOut_3 <= lengths_47;
            end else if (8'h2e == characterIndex) begin
              lengthsOut_3 <= lengths_46;
            end else if (8'h2d == characterIndex) begin
              lengthsOut_3 <= lengths_45;
            end else if (8'h2c == characterIndex) begin
              lengthsOut_3 <= lengths_44;
            end else if (8'h2b == characterIndex) begin
              lengthsOut_3 <= lengths_43;
            end else if (8'h2a == characterIndex) begin
              lengthsOut_3 <= lengths_42;
            end else if (8'h29 == characterIndex) begin
              lengthsOut_3 <= lengths_41;
            end else if (8'h28 == characterIndex) begin
              lengthsOut_3 <= lengths_40;
            end else if (8'h27 == characterIndex) begin
              lengthsOut_3 <= lengths_39;
            end else if (8'h26 == characterIndex) begin
              lengthsOut_3 <= lengths_38;
            end else if (8'h25 == characterIndex) begin
              lengthsOut_3 <= lengths_37;
            end else if (8'h24 == characterIndex) begin
              lengthsOut_3 <= lengths_36;
            end else if (8'h23 == characterIndex) begin
              lengthsOut_3 <= lengths_35;
            end else if (8'h22 == characterIndex) begin
              lengthsOut_3 <= lengths_34;
            end else if (8'h21 == characterIndex) begin
              lengthsOut_3 <= lengths_33;
            end else if (8'h20 == characterIndex) begin
              lengthsOut_3 <= lengths_32;
            end else if (8'h1f == characterIndex) begin
              lengthsOut_3 <= lengths_31;
            end else if (8'h1e == characterIndex) begin
              lengthsOut_3 <= lengths_30;
            end else if (8'h1d == characterIndex) begin
              lengthsOut_3 <= lengths_29;
            end else if (8'h1c == characterIndex) begin
              lengthsOut_3 <= lengths_28;
            end else if (8'h1b == characterIndex) begin
              lengthsOut_3 <= lengths_27;
            end else if (8'h1a == characterIndex) begin
              lengthsOut_3 <= lengths_26;
            end else if (8'h19 == characterIndex) begin
              lengthsOut_3 <= lengths_25;
            end else if (8'h18 == characterIndex) begin
              lengthsOut_3 <= lengths_24;
            end else if (8'h17 == characterIndex) begin
              lengthsOut_3 <= lengths_23;
            end else if (8'h16 == characterIndex) begin
              lengthsOut_3 <= lengths_22;
            end else if (8'h15 == characterIndex) begin
              lengthsOut_3 <= lengths_21;
            end else if (8'h14 == characterIndex) begin
              lengthsOut_3 <= lengths_20;
            end else if (8'h13 == characterIndex) begin
              lengthsOut_3 <= lengths_19;
            end else if (8'h12 == characterIndex) begin
              lengthsOut_3 <= lengths_18;
            end else if (8'h11 == characterIndex) begin
              lengthsOut_3 <= lengths_17;
            end else if (8'h10 == characterIndex) begin
              lengthsOut_3 <= lengths_16;
            end else if (8'hf == characterIndex) begin
              lengthsOut_3 <= lengths_15;
            end else if (8'he == characterIndex) begin
              lengthsOut_3 <= lengths_14;
            end else if (8'hd == characterIndex) begin
              lengthsOut_3 <= lengths_13;
            end else if (8'hc == characterIndex) begin
              lengthsOut_3 <= lengths_12;
            end else if (8'hb == characterIndex) begin
              lengthsOut_3 <= lengths_11;
            end else if (8'ha == characterIndex) begin
              lengthsOut_3 <= lengths_10;
            end else if (8'h9 == characterIndex) begin
              lengthsOut_3 <= lengths_9;
            end else if (8'h8 == characterIndex) begin
              lengthsOut_3 <= lengths_8;
            end else if (8'h7 == characterIndex) begin
              lengthsOut_3 <= lengths_7;
            end else if (8'h6 == characterIndex) begin
              lengthsOut_3 <= lengths_6;
            end else if (8'h5 == characterIndex) begin
              lengthsOut_3 <= lengths_5;
            end else if (8'h4 == characterIndex) begin
              lengthsOut_3 <= lengths_4;
            end else if (8'h3 == characterIndex) begin
              lengthsOut_3 <= lengths_3;
            end else if (8'h2 == characterIndex) begin
              lengthsOut_3 <= lengths_2;
            end else if (8'h1 == characterIndex) begin
              lengthsOut_3 <= lengths_1;
            end else begin
              lengthsOut_3 <= lengths_0;
            end
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h4 == characterIndex) begin
              lengthsOut_4 <= _T_69;
            end
          end else if (8'h4 == characterIndex) begin
            lengthsOut_4 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h5 == characterIndex) begin
              lengthsOut_5 <= _T_69;
            end
          end else if (8'h5 == characterIndex) begin
            lengthsOut_5 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h6 == characterIndex) begin
              lengthsOut_6 <= _T_69;
            end
          end else if (8'h6 == characterIndex) begin
            lengthsOut_6 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h7 == characterIndex) begin
              lengthsOut_7 <= _T_69;
            end
          end else if (8'h7 == characterIndex) begin
            lengthsOut_7 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h8 == characterIndex) begin
              lengthsOut_8 <= _T_69;
            end
          end else if (8'h8 == characterIndex) begin
            lengthsOut_8 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h9 == characterIndex) begin
              lengthsOut_9 <= _T_69;
            end
          end else if (8'h9 == characterIndex) begin
            lengthsOut_9 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha == characterIndex) begin
              lengthsOut_10 <= _T_69;
            end
          end else if (8'ha == characterIndex) begin
            lengthsOut_10 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb == characterIndex) begin
              lengthsOut_11 <= _T_69;
            end
          end else if (8'hb == characterIndex) begin
            lengthsOut_11 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc == characterIndex) begin
              lengthsOut_12 <= _T_69;
            end
          end else if (8'hc == characterIndex) begin
            lengthsOut_12 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd == characterIndex) begin
              lengthsOut_13 <= _T_69;
            end
          end else if (8'hd == characterIndex) begin
            lengthsOut_13 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he == characterIndex) begin
              lengthsOut_14 <= _T_69;
            end
          end else if (8'he == characterIndex) begin
            lengthsOut_14 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf == characterIndex) begin
              lengthsOut_15 <= _T_69;
            end
          end else if (8'hf == characterIndex) begin
            lengthsOut_15 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h10 == characterIndex) begin
              lengthsOut_16 <= _T_69;
            end
          end else if (8'h10 == characterIndex) begin
            lengthsOut_16 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h11 == characterIndex) begin
              lengthsOut_17 <= _T_69;
            end
          end else if (8'h11 == characterIndex) begin
            lengthsOut_17 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h12 == characterIndex) begin
              lengthsOut_18 <= _T_69;
            end
          end else if (8'h12 == characterIndex) begin
            lengthsOut_18 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h13 == characterIndex) begin
              lengthsOut_19 <= _T_69;
            end
          end else if (8'h13 == characterIndex) begin
            lengthsOut_19 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h14 == characterIndex) begin
              lengthsOut_20 <= _T_69;
            end
          end else if (8'h14 == characterIndex) begin
            lengthsOut_20 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h15 == characterIndex) begin
              lengthsOut_21 <= _T_69;
            end
          end else if (8'h15 == characterIndex) begin
            lengthsOut_21 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h16 == characterIndex) begin
              lengthsOut_22 <= _T_69;
            end
          end else if (8'h16 == characterIndex) begin
            lengthsOut_22 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h17 == characterIndex) begin
              lengthsOut_23 <= _T_69;
            end
          end else if (8'h17 == characterIndex) begin
            lengthsOut_23 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h18 == characterIndex) begin
              lengthsOut_24 <= _T_69;
            end
          end else if (8'h18 == characterIndex) begin
            lengthsOut_24 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h19 == characterIndex) begin
              lengthsOut_25 <= _T_69;
            end
          end else if (8'h19 == characterIndex) begin
            lengthsOut_25 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h1a == characterIndex) begin
              lengthsOut_26 <= _T_69;
            end
          end else if (8'h1a == characterIndex) begin
            lengthsOut_26 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h1b == characterIndex) begin
              lengthsOut_27 <= _T_69;
            end
          end else if (8'h1b == characterIndex) begin
            lengthsOut_27 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h1c == characterIndex) begin
              lengthsOut_28 <= _T_69;
            end
          end else if (8'h1c == characterIndex) begin
            lengthsOut_28 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h1d == characterIndex) begin
              lengthsOut_29 <= _T_69;
            end
          end else if (8'h1d == characterIndex) begin
            lengthsOut_29 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h1e == characterIndex) begin
              lengthsOut_30 <= _T_69;
            end
          end else if (8'h1e == characterIndex) begin
            lengthsOut_30 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h1f == characterIndex) begin
              lengthsOut_31 <= _T_69;
            end
          end else if (8'h1f == characterIndex) begin
            lengthsOut_31 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h20 == characterIndex) begin
              lengthsOut_32 <= _T_69;
            end
          end else if (8'h20 == characterIndex) begin
            lengthsOut_32 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h21 == characterIndex) begin
              lengthsOut_33 <= _T_69;
            end
          end else if (8'h21 == characterIndex) begin
            lengthsOut_33 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h22 == characterIndex) begin
              lengthsOut_34 <= _T_69;
            end
          end else if (8'h22 == characterIndex) begin
            lengthsOut_34 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h23 == characterIndex) begin
              lengthsOut_35 <= _T_69;
            end
          end else if (8'h23 == characterIndex) begin
            lengthsOut_35 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h24 == characterIndex) begin
              lengthsOut_36 <= _T_69;
            end
          end else if (8'h24 == characterIndex) begin
            lengthsOut_36 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h25 == characterIndex) begin
              lengthsOut_37 <= _T_69;
            end
          end else if (8'h25 == characterIndex) begin
            lengthsOut_37 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h26 == characterIndex) begin
              lengthsOut_38 <= _T_69;
            end
          end else if (8'h26 == characterIndex) begin
            lengthsOut_38 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h27 == characterIndex) begin
              lengthsOut_39 <= _T_69;
            end
          end else if (8'h27 == characterIndex) begin
            lengthsOut_39 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h28 == characterIndex) begin
              lengthsOut_40 <= _T_69;
            end
          end else if (8'h28 == characterIndex) begin
            lengthsOut_40 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h29 == characterIndex) begin
              lengthsOut_41 <= _T_69;
            end
          end else if (8'h29 == characterIndex) begin
            lengthsOut_41 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h2a == characterIndex) begin
              lengthsOut_42 <= _T_69;
            end
          end else if (8'h2a == characterIndex) begin
            lengthsOut_42 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h2b == characterIndex) begin
              lengthsOut_43 <= _T_69;
            end
          end else if (8'h2b == characterIndex) begin
            lengthsOut_43 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h2c == characterIndex) begin
              lengthsOut_44 <= _T_69;
            end
          end else if (8'h2c == characterIndex) begin
            lengthsOut_44 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h2d == characterIndex) begin
              lengthsOut_45 <= _T_69;
            end
          end else if (8'h2d == characterIndex) begin
            lengthsOut_45 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h2e == characterIndex) begin
              lengthsOut_46 <= _T_69;
            end
          end else if (8'h2e == characterIndex) begin
            lengthsOut_46 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h2f == characterIndex) begin
              lengthsOut_47 <= _T_69;
            end
          end else if (8'h2f == characterIndex) begin
            lengthsOut_47 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h30 == characterIndex) begin
              lengthsOut_48 <= _T_69;
            end
          end else if (8'h30 == characterIndex) begin
            lengthsOut_48 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h31 == characterIndex) begin
              lengthsOut_49 <= _T_69;
            end
          end else if (8'h31 == characterIndex) begin
            lengthsOut_49 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h32 == characterIndex) begin
              lengthsOut_50 <= _T_69;
            end
          end else if (8'h32 == characterIndex) begin
            lengthsOut_50 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h33 == characterIndex) begin
              lengthsOut_51 <= _T_69;
            end
          end else if (8'h33 == characterIndex) begin
            lengthsOut_51 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h34 == characterIndex) begin
              lengthsOut_52 <= _T_69;
            end
          end else if (8'h34 == characterIndex) begin
            lengthsOut_52 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h35 == characterIndex) begin
              lengthsOut_53 <= _T_69;
            end
          end else if (8'h35 == characterIndex) begin
            lengthsOut_53 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h36 == characterIndex) begin
              lengthsOut_54 <= _T_69;
            end
          end else if (8'h36 == characterIndex) begin
            lengthsOut_54 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h37 == characterIndex) begin
              lengthsOut_55 <= _T_69;
            end
          end else if (8'h37 == characterIndex) begin
            lengthsOut_55 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h38 == characterIndex) begin
              lengthsOut_56 <= _T_69;
            end
          end else if (8'h38 == characterIndex) begin
            lengthsOut_56 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h39 == characterIndex) begin
              lengthsOut_57 <= _T_69;
            end
          end else if (8'h39 == characterIndex) begin
            lengthsOut_57 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h3a == characterIndex) begin
              lengthsOut_58 <= _T_69;
            end
          end else if (8'h3a == characterIndex) begin
            lengthsOut_58 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h3b == characterIndex) begin
              lengthsOut_59 <= _T_69;
            end
          end else if (8'h3b == characterIndex) begin
            lengthsOut_59 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h3c == characterIndex) begin
              lengthsOut_60 <= _T_69;
            end
          end else if (8'h3c == characterIndex) begin
            lengthsOut_60 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h3d == characterIndex) begin
              lengthsOut_61 <= _T_69;
            end
          end else if (8'h3d == characterIndex) begin
            lengthsOut_61 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h3e == characterIndex) begin
              lengthsOut_62 <= _T_69;
            end
          end else if (8'h3e == characterIndex) begin
            lengthsOut_62 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h3f == characterIndex) begin
              lengthsOut_63 <= _T_69;
            end
          end else if (8'h3f == characterIndex) begin
            lengthsOut_63 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h40 == characterIndex) begin
              lengthsOut_64 <= _T_69;
            end
          end else if (8'h40 == characterIndex) begin
            lengthsOut_64 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h41 == characterIndex) begin
              lengthsOut_65 <= _T_69;
            end
          end else if (8'h41 == characterIndex) begin
            lengthsOut_65 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h42 == characterIndex) begin
              lengthsOut_66 <= _T_69;
            end
          end else if (8'h42 == characterIndex) begin
            lengthsOut_66 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h43 == characterIndex) begin
              lengthsOut_67 <= _T_69;
            end
          end else if (8'h43 == characterIndex) begin
            lengthsOut_67 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h44 == characterIndex) begin
              lengthsOut_68 <= _T_69;
            end
          end else if (8'h44 == characterIndex) begin
            lengthsOut_68 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h45 == characterIndex) begin
              lengthsOut_69 <= _T_69;
            end
          end else if (8'h45 == characterIndex) begin
            lengthsOut_69 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h46 == characterIndex) begin
              lengthsOut_70 <= _T_69;
            end
          end else if (8'h46 == characterIndex) begin
            lengthsOut_70 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h47 == characterIndex) begin
              lengthsOut_71 <= _T_69;
            end
          end else if (8'h47 == characterIndex) begin
            lengthsOut_71 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h48 == characterIndex) begin
              lengthsOut_72 <= _T_69;
            end
          end else if (8'h48 == characterIndex) begin
            lengthsOut_72 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h49 == characterIndex) begin
              lengthsOut_73 <= _T_69;
            end
          end else if (8'h49 == characterIndex) begin
            lengthsOut_73 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h4a == characterIndex) begin
              lengthsOut_74 <= _T_69;
            end
          end else if (8'h4a == characterIndex) begin
            lengthsOut_74 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h4b == characterIndex) begin
              lengthsOut_75 <= _T_69;
            end
          end else if (8'h4b == characterIndex) begin
            lengthsOut_75 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h4c == characterIndex) begin
              lengthsOut_76 <= _T_69;
            end
          end else if (8'h4c == characterIndex) begin
            lengthsOut_76 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h4d == characterIndex) begin
              lengthsOut_77 <= _T_69;
            end
          end else if (8'h4d == characterIndex) begin
            lengthsOut_77 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h4e == characterIndex) begin
              lengthsOut_78 <= _T_69;
            end
          end else if (8'h4e == characterIndex) begin
            lengthsOut_78 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h4f == characterIndex) begin
              lengthsOut_79 <= _T_69;
            end
          end else if (8'h4f == characterIndex) begin
            lengthsOut_79 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h50 == characterIndex) begin
              lengthsOut_80 <= _T_69;
            end
          end else if (8'h50 == characterIndex) begin
            lengthsOut_80 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h51 == characterIndex) begin
              lengthsOut_81 <= _T_69;
            end
          end else if (8'h51 == characterIndex) begin
            lengthsOut_81 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h52 == characterIndex) begin
              lengthsOut_82 <= _T_69;
            end
          end else if (8'h52 == characterIndex) begin
            lengthsOut_82 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h53 == characterIndex) begin
              lengthsOut_83 <= _T_69;
            end
          end else if (8'h53 == characterIndex) begin
            lengthsOut_83 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h54 == characterIndex) begin
              lengthsOut_84 <= _T_69;
            end
          end else if (8'h54 == characterIndex) begin
            lengthsOut_84 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h55 == characterIndex) begin
              lengthsOut_85 <= _T_69;
            end
          end else if (8'h55 == characterIndex) begin
            lengthsOut_85 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h56 == characterIndex) begin
              lengthsOut_86 <= _T_69;
            end
          end else if (8'h56 == characterIndex) begin
            lengthsOut_86 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h57 == characterIndex) begin
              lengthsOut_87 <= _T_69;
            end
          end else if (8'h57 == characterIndex) begin
            lengthsOut_87 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h58 == characterIndex) begin
              lengthsOut_88 <= _T_69;
            end
          end else if (8'h58 == characterIndex) begin
            lengthsOut_88 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h59 == characterIndex) begin
              lengthsOut_89 <= _T_69;
            end
          end else if (8'h59 == characterIndex) begin
            lengthsOut_89 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h5a == characterIndex) begin
              lengthsOut_90 <= _T_69;
            end
          end else if (8'h5a == characterIndex) begin
            lengthsOut_90 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h5b == characterIndex) begin
              lengthsOut_91 <= _T_69;
            end
          end else if (8'h5b == characterIndex) begin
            lengthsOut_91 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h5c == characterIndex) begin
              lengthsOut_92 <= _T_69;
            end
          end else if (8'h5c == characterIndex) begin
            lengthsOut_92 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h5d == characterIndex) begin
              lengthsOut_93 <= _T_69;
            end
          end else if (8'h5d == characterIndex) begin
            lengthsOut_93 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h5e == characterIndex) begin
              lengthsOut_94 <= _T_69;
            end
          end else if (8'h5e == characterIndex) begin
            lengthsOut_94 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h5f == characterIndex) begin
              lengthsOut_95 <= _T_69;
            end
          end else if (8'h5f == characterIndex) begin
            lengthsOut_95 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h60 == characterIndex) begin
              lengthsOut_96 <= _T_69;
            end
          end else if (8'h60 == characterIndex) begin
            lengthsOut_96 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h61 == characterIndex) begin
              lengthsOut_97 <= _T_69;
            end
          end else if (8'h61 == characterIndex) begin
            lengthsOut_97 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h62 == characterIndex) begin
              lengthsOut_98 <= _T_69;
            end
          end else if (8'h62 == characterIndex) begin
            lengthsOut_98 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h63 == characterIndex) begin
              lengthsOut_99 <= _T_69;
            end
          end else if (8'h63 == characterIndex) begin
            lengthsOut_99 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h64 == characterIndex) begin
              lengthsOut_100 <= _T_69;
            end
          end else if (8'h64 == characterIndex) begin
            lengthsOut_100 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h65 == characterIndex) begin
              lengthsOut_101 <= _T_69;
            end
          end else if (8'h65 == characterIndex) begin
            lengthsOut_101 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h66 == characterIndex) begin
              lengthsOut_102 <= _T_69;
            end
          end else if (8'h66 == characterIndex) begin
            lengthsOut_102 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h67 == characterIndex) begin
              lengthsOut_103 <= _T_69;
            end
          end else if (8'h67 == characterIndex) begin
            lengthsOut_103 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h68 == characterIndex) begin
              lengthsOut_104 <= _T_69;
            end
          end else if (8'h68 == characterIndex) begin
            lengthsOut_104 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h69 == characterIndex) begin
              lengthsOut_105 <= _T_69;
            end
          end else if (8'h69 == characterIndex) begin
            lengthsOut_105 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h6a == characterIndex) begin
              lengthsOut_106 <= _T_69;
            end
          end else if (8'h6a == characterIndex) begin
            lengthsOut_106 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h6b == characterIndex) begin
              lengthsOut_107 <= _T_69;
            end
          end else if (8'h6b == characterIndex) begin
            lengthsOut_107 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h6c == characterIndex) begin
              lengthsOut_108 <= _T_69;
            end
          end else if (8'h6c == characterIndex) begin
            lengthsOut_108 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h6d == characterIndex) begin
              lengthsOut_109 <= _T_69;
            end
          end else if (8'h6d == characterIndex) begin
            lengthsOut_109 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h6e == characterIndex) begin
              lengthsOut_110 <= _T_69;
            end
          end else if (8'h6e == characterIndex) begin
            lengthsOut_110 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h6f == characterIndex) begin
              lengthsOut_111 <= _T_69;
            end
          end else if (8'h6f == characterIndex) begin
            lengthsOut_111 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h70 == characterIndex) begin
              lengthsOut_112 <= _T_69;
            end
          end else if (8'h70 == characterIndex) begin
            lengthsOut_112 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h71 == characterIndex) begin
              lengthsOut_113 <= _T_69;
            end
          end else if (8'h71 == characterIndex) begin
            lengthsOut_113 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h72 == characterIndex) begin
              lengthsOut_114 <= _T_69;
            end
          end else if (8'h72 == characterIndex) begin
            lengthsOut_114 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h73 == characterIndex) begin
              lengthsOut_115 <= _T_69;
            end
          end else if (8'h73 == characterIndex) begin
            lengthsOut_115 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h74 == characterIndex) begin
              lengthsOut_116 <= _T_69;
            end
          end else if (8'h74 == characterIndex) begin
            lengthsOut_116 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h75 == characterIndex) begin
              lengthsOut_117 <= _T_69;
            end
          end else if (8'h75 == characterIndex) begin
            lengthsOut_117 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h76 == characterIndex) begin
              lengthsOut_118 <= _T_69;
            end
          end else if (8'h76 == characterIndex) begin
            lengthsOut_118 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h77 == characterIndex) begin
              lengthsOut_119 <= _T_69;
            end
          end else if (8'h77 == characterIndex) begin
            lengthsOut_119 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h78 == characterIndex) begin
              lengthsOut_120 <= _T_69;
            end
          end else if (8'h78 == characterIndex) begin
            lengthsOut_120 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h79 == characterIndex) begin
              lengthsOut_121 <= _T_69;
            end
          end else if (8'h79 == characterIndex) begin
            lengthsOut_121 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h7a == characterIndex) begin
              lengthsOut_122 <= _T_69;
            end
          end else if (8'h7a == characterIndex) begin
            lengthsOut_122 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h7b == characterIndex) begin
              lengthsOut_123 <= _T_69;
            end
          end else if (8'h7b == characterIndex) begin
            lengthsOut_123 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h7c == characterIndex) begin
              lengthsOut_124 <= _T_69;
            end
          end else if (8'h7c == characterIndex) begin
            lengthsOut_124 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h7d == characterIndex) begin
              lengthsOut_125 <= _T_69;
            end
          end else if (8'h7d == characterIndex) begin
            lengthsOut_125 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h7e == characterIndex) begin
              lengthsOut_126 <= _T_69;
            end
          end else if (8'h7e == characterIndex) begin
            lengthsOut_126 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h7f == characterIndex) begin
              lengthsOut_127 <= _T_69;
            end
          end else if (8'h7f == characterIndex) begin
            lengthsOut_127 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h80 == characterIndex) begin
              lengthsOut_128 <= _T_69;
            end
          end else if (8'h80 == characterIndex) begin
            lengthsOut_128 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h81 == characterIndex) begin
              lengthsOut_129 <= _T_69;
            end
          end else if (8'h81 == characterIndex) begin
            lengthsOut_129 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h82 == characterIndex) begin
              lengthsOut_130 <= _T_69;
            end
          end else if (8'h82 == characterIndex) begin
            lengthsOut_130 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h83 == characterIndex) begin
              lengthsOut_131 <= _T_69;
            end
          end else if (8'h83 == characterIndex) begin
            lengthsOut_131 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h84 == characterIndex) begin
              lengthsOut_132 <= _T_69;
            end
          end else if (8'h84 == characterIndex) begin
            lengthsOut_132 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h85 == characterIndex) begin
              lengthsOut_133 <= _T_69;
            end
          end else if (8'h85 == characterIndex) begin
            lengthsOut_133 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h86 == characterIndex) begin
              lengthsOut_134 <= _T_69;
            end
          end else if (8'h86 == characterIndex) begin
            lengthsOut_134 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h87 == characterIndex) begin
              lengthsOut_135 <= _T_69;
            end
          end else if (8'h87 == characterIndex) begin
            lengthsOut_135 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h88 == characterIndex) begin
              lengthsOut_136 <= _T_69;
            end
          end else if (8'h88 == characterIndex) begin
            lengthsOut_136 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h89 == characterIndex) begin
              lengthsOut_137 <= _T_69;
            end
          end else if (8'h89 == characterIndex) begin
            lengthsOut_137 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h8a == characterIndex) begin
              lengthsOut_138 <= _T_69;
            end
          end else if (8'h8a == characterIndex) begin
            lengthsOut_138 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h8b == characterIndex) begin
              lengthsOut_139 <= _T_69;
            end
          end else if (8'h8b == characterIndex) begin
            lengthsOut_139 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h8c == characterIndex) begin
              lengthsOut_140 <= _T_69;
            end
          end else if (8'h8c == characterIndex) begin
            lengthsOut_140 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h8d == characterIndex) begin
              lengthsOut_141 <= _T_69;
            end
          end else if (8'h8d == characterIndex) begin
            lengthsOut_141 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h8e == characterIndex) begin
              lengthsOut_142 <= _T_69;
            end
          end else if (8'h8e == characterIndex) begin
            lengthsOut_142 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h8f == characterIndex) begin
              lengthsOut_143 <= _T_69;
            end
          end else if (8'h8f == characterIndex) begin
            lengthsOut_143 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h90 == characterIndex) begin
              lengthsOut_144 <= _T_69;
            end
          end else if (8'h90 == characterIndex) begin
            lengthsOut_144 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h91 == characterIndex) begin
              lengthsOut_145 <= _T_69;
            end
          end else if (8'h91 == characterIndex) begin
            lengthsOut_145 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h92 == characterIndex) begin
              lengthsOut_146 <= _T_69;
            end
          end else if (8'h92 == characterIndex) begin
            lengthsOut_146 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h93 == characterIndex) begin
              lengthsOut_147 <= _T_69;
            end
          end else if (8'h93 == characterIndex) begin
            lengthsOut_147 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h94 == characterIndex) begin
              lengthsOut_148 <= _T_69;
            end
          end else if (8'h94 == characterIndex) begin
            lengthsOut_148 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h95 == characterIndex) begin
              lengthsOut_149 <= _T_69;
            end
          end else if (8'h95 == characterIndex) begin
            lengthsOut_149 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h96 == characterIndex) begin
              lengthsOut_150 <= _T_69;
            end
          end else if (8'h96 == characterIndex) begin
            lengthsOut_150 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h97 == characterIndex) begin
              lengthsOut_151 <= _T_69;
            end
          end else if (8'h97 == characterIndex) begin
            lengthsOut_151 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h98 == characterIndex) begin
              lengthsOut_152 <= _T_69;
            end
          end else if (8'h98 == characterIndex) begin
            lengthsOut_152 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h99 == characterIndex) begin
              lengthsOut_153 <= _T_69;
            end
          end else if (8'h99 == characterIndex) begin
            lengthsOut_153 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h9a == characterIndex) begin
              lengthsOut_154 <= _T_69;
            end
          end else if (8'h9a == characterIndex) begin
            lengthsOut_154 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h9b == characterIndex) begin
              lengthsOut_155 <= _T_69;
            end
          end else if (8'h9b == characterIndex) begin
            lengthsOut_155 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h9c == characterIndex) begin
              lengthsOut_156 <= _T_69;
            end
          end else if (8'h9c == characterIndex) begin
            lengthsOut_156 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h9d == characterIndex) begin
              lengthsOut_157 <= _T_69;
            end
          end else if (8'h9d == characterIndex) begin
            lengthsOut_157 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h9e == characterIndex) begin
              lengthsOut_158 <= _T_69;
            end
          end else if (8'h9e == characterIndex) begin
            lengthsOut_158 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'h9f == characterIndex) begin
              lengthsOut_159 <= _T_69;
            end
          end else if (8'h9f == characterIndex) begin
            lengthsOut_159 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha0 == characterIndex) begin
              lengthsOut_160 <= _T_69;
            end
          end else if (8'ha0 == characterIndex) begin
            lengthsOut_160 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha1 == characterIndex) begin
              lengthsOut_161 <= _T_69;
            end
          end else if (8'ha1 == characterIndex) begin
            lengthsOut_161 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha2 == characterIndex) begin
              lengthsOut_162 <= _T_69;
            end
          end else if (8'ha2 == characterIndex) begin
            lengthsOut_162 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha3 == characterIndex) begin
              lengthsOut_163 <= _T_69;
            end
          end else if (8'ha3 == characterIndex) begin
            lengthsOut_163 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha4 == characterIndex) begin
              lengthsOut_164 <= _T_69;
            end
          end else if (8'ha4 == characterIndex) begin
            lengthsOut_164 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha5 == characterIndex) begin
              lengthsOut_165 <= _T_69;
            end
          end else if (8'ha5 == characterIndex) begin
            lengthsOut_165 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha6 == characterIndex) begin
              lengthsOut_166 <= _T_69;
            end
          end else if (8'ha6 == characterIndex) begin
            lengthsOut_166 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha7 == characterIndex) begin
              lengthsOut_167 <= _T_69;
            end
          end else if (8'ha7 == characterIndex) begin
            lengthsOut_167 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha8 == characterIndex) begin
              lengthsOut_168 <= _T_69;
            end
          end else if (8'ha8 == characterIndex) begin
            lengthsOut_168 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'ha9 == characterIndex) begin
              lengthsOut_169 <= _T_69;
            end
          end else if (8'ha9 == characterIndex) begin
            lengthsOut_169 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'haa == characterIndex) begin
              lengthsOut_170 <= _T_69;
            end
          end else if (8'haa == characterIndex) begin
            lengthsOut_170 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hab == characterIndex) begin
              lengthsOut_171 <= _T_69;
            end
          end else if (8'hab == characterIndex) begin
            lengthsOut_171 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hac == characterIndex) begin
              lengthsOut_172 <= _T_69;
            end
          end else if (8'hac == characterIndex) begin
            lengthsOut_172 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'had == characterIndex) begin
              lengthsOut_173 <= _T_69;
            end
          end else if (8'had == characterIndex) begin
            lengthsOut_173 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hae == characterIndex) begin
              lengthsOut_174 <= _T_69;
            end
          end else if (8'hae == characterIndex) begin
            lengthsOut_174 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'haf == characterIndex) begin
              lengthsOut_175 <= _T_69;
            end
          end else if (8'haf == characterIndex) begin
            lengthsOut_175 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb0 == characterIndex) begin
              lengthsOut_176 <= _T_69;
            end
          end else if (8'hb0 == characterIndex) begin
            lengthsOut_176 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb1 == characterIndex) begin
              lengthsOut_177 <= _T_69;
            end
          end else if (8'hb1 == characterIndex) begin
            lengthsOut_177 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb2 == characterIndex) begin
              lengthsOut_178 <= _T_69;
            end
          end else if (8'hb2 == characterIndex) begin
            lengthsOut_178 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb3 == characterIndex) begin
              lengthsOut_179 <= _T_69;
            end
          end else if (8'hb3 == characterIndex) begin
            lengthsOut_179 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb4 == characterIndex) begin
              lengthsOut_180 <= _T_69;
            end
          end else if (8'hb4 == characterIndex) begin
            lengthsOut_180 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb5 == characterIndex) begin
              lengthsOut_181 <= _T_69;
            end
          end else if (8'hb5 == characterIndex) begin
            lengthsOut_181 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb6 == characterIndex) begin
              lengthsOut_182 <= _T_69;
            end
          end else if (8'hb6 == characterIndex) begin
            lengthsOut_182 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb7 == characterIndex) begin
              lengthsOut_183 <= _T_69;
            end
          end else if (8'hb7 == characterIndex) begin
            lengthsOut_183 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb8 == characterIndex) begin
              lengthsOut_184 <= _T_69;
            end
          end else if (8'hb8 == characterIndex) begin
            lengthsOut_184 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hb9 == characterIndex) begin
              lengthsOut_185 <= _T_69;
            end
          end else if (8'hb9 == characterIndex) begin
            lengthsOut_185 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hba == characterIndex) begin
              lengthsOut_186 <= _T_69;
            end
          end else if (8'hba == characterIndex) begin
            lengthsOut_186 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hbb == characterIndex) begin
              lengthsOut_187 <= _T_69;
            end
          end else if (8'hbb == characterIndex) begin
            lengthsOut_187 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hbc == characterIndex) begin
              lengthsOut_188 <= _T_69;
            end
          end else if (8'hbc == characterIndex) begin
            lengthsOut_188 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hbd == characterIndex) begin
              lengthsOut_189 <= _T_69;
            end
          end else if (8'hbd == characterIndex) begin
            lengthsOut_189 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hbe == characterIndex) begin
              lengthsOut_190 <= _T_69;
            end
          end else if (8'hbe == characterIndex) begin
            lengthsOut_190 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hbf == characterIndex) begin
              lengthsOut_191 <= _T_69;
            end
          end else if (8'hbf == characterIndex) begin
            lengthsOut_191 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc0 == characterIndex) begin
              lengthsOut_192 <= _T_69;
            end
          end else if (8'hc0 == characterIndex) begin
            lengthsOut_192 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc1 == characterIndex) begin
              lengthsOut_193 <= _T_69;
            end
          end else if (8'hc1 == characterIndex) begin
            lengthsOut_193 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc2 == characterIndex) begin
              lengthsOut_194 <= _T_69;
            end
          end else if (8'hc2 == characterIndex) begin
            lengthsOut_194 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc3 == characterIndex) begin
              lengthsOut_195 <= _T_69;
            end
          end else if (8'hc3 == characterIndex) begin
            lengthsOut_195 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc4 == characterIndex) begin
              lengthsOut_196 <= _T_69;
            end
          end else if (8'hc4 == characterIndex) begin
            lengthsOut_196 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc5 == characterIndex) begin
              lengthsOut_197 <= _T_69;
            end
          end else if (8'hc5 == characterIndex) begin
            lengthsOut_197 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc6 == characterIndex) begin
              lengthsOut_198 <= _T_69;
            end
          end else if (8'hc6 == characterIndex) begin
            lengthsOut_198 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc7 == characterIndex) begin
              lengthsOut_199 <= _T_69;
            end
          end else if (8'hc7 == characterIndex) begin
            lengthsOut_199 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc8 == characterIndex) begin
              lengthsOut_200 <= _T_69;
            end
          end else if (8'hc8 == characterIndex) begin
            lengthsOut_200 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hc9 == characterIndex) begin
              lengthsOut_201 <= _T_69;
            end
          end else if (8'hc9 == characterIndex) begin
            lengthsOut_201 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hca == characterIndex) begin
              lengthsOut_202 <= _T_69;
            end
          end else if (8'hca == characterIndex) begin
            lengthsOut_202 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hcb == characterIndex) begin
              lengthsOut_203 <= _T_69;
            end
          end else if (8'hcb == characterIndex) begin
            lengthsOut_203 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hcc == characterIndex) begin
              lengthsOut_204 <= _T_69;
            end
          end else if (8'hcc == characterIndex) begin
            lengthsOut_204 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hcd == characterIndex) begin
              lengthsOut_205 <= _T_69;
            end
          end else if (8'hcd == characterIndex) begin
            lengthsOut_205 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hce == characterIndex) begin
              lengthsOut_206 <= _T_69;
            end
          end else if (8'hce == characterIndex) begin
            lengthsOut_206 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hcf == characterIndex) begin
              lengthsOut_207 <= _T_69;
            end
          end else if (8'hcf == characterIndex) begin
            lengthsOut_207 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd0 == characterIndex) begin
              lengthsOut_208 <= _T_69;
            end
          end else if (8'hd0 == characterIndex) begin
            lengthsOut_208 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd1 == characterIndex) begin
              lengthsOut_209 <= _T_69;
            end
          end else if (8'hd1 == characterIndex) begin
            lengthsOut_209 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd2 == characterIndex) begin
              lengthsOut_210 <= _T_69;
            end
          end else if (8'hd2 == characterIndex) begin
            lengthsOut_210 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd3 == characterIndex) begin
              lengthsOut_211 <= _T_69;
            end
          end else if (8'hd3 == characterIndex) begin
            lengthsOut_211 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd4 == characterIndex) begin
              lengthsOut_212 <= _T_69;
            end
          end else if (8'hd4 == characterIndex) begin
            lengthsOut_212 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd5 == characterIndex) begin
              lengthsOut_213 <= _T_69;
            end
          end else if (8'hd5 == characterIndex) begin
            lengthsOut_213 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd6 == characterIndex) begin
              lengthsOut_214 <= _T_69;
            end
          end else if (8'hd6 == characterIndex) begin
            lengthsOut_214 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd7 == characterIndex) begin
              lengthsOut_215 <= _T_69;
            end
          end else if (8'hd7 == characterIndex) begin
            lengthsOut_215 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd8 == characterIndex) begin
              lengthsOut_216 <= _T_69;
            end
          end else if (8'hd8 == characterIndex) begin
            lengthsOut_216 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hd9 == characterIndex) begin
              lengthsOut_217 <= _T_69;
            end
          end else if (8'hd9 == characterIndex) begin
            lengthsOut_217 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hda == characterIndex) begin
              lengthsOut_218 <= _T_69;
            end
          end else if (8'hda == characterIndex) begin
            lengthsOut_218 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hdb == characterIndex) begin
              lengthsOut_219 <= _T_69;
            end
          end else if (8'hdb == characterIndex) begin
            lengthsOut_219 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hdc == characterIndex) begin
              lengthsOut_220 <= _T_69;
            end
          end else if (8'hdc == characterIndex) begin
            lengthsOut_220 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hdd == characterIndex) begin
              lengthsOut_221 <= _T_69;
            end
          end else if (8'hdd == characterIndex) begin
            lengthsOut_221 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hde == characterIndex) begin
              lengthsOut_222 <= _T_69;
            end
          end else if (8'hde == characterIndex) begin
            lengthsOut_222 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hdf == characterIndex) begin
              lengthsOut_223 <= _T_69;
            end
          end else if (8'hdf == characterIndex) begin
            lengthsOut_223 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he0 == characterIndex) begin
              lengthsOut_224 <= _T_69;
            end
          end else if (8'he0 == characterIndex) begin
            lengthsOut_224 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he1 == characterIndex) begin
              lengthsOut_225 <= _T_69;
            end
          end else if (8'he1 == characterIndex) begin
            lengthsOut_225 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he2 == characterIndex) begin
              lengthsOut_226 <= _T_69;
            end
          end else if (8'he2 == characterIndex) begin
            lengthsOut_226 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he3 == characterIndex) begin
              lengthsOut_227 <= _T_69;
            end
          end else if (8'he3 == characterIndex) begin
            lengthsOut_227 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he4 == characterIndex) begin
              lengthsOut_228 <= _T_69;
            end
          end else if (8'he4 == characterIndex) begin
            lengthsOut_228 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he5 == characterIndex) begin
              lengthsOut_229 <= _T_69;
            end
          end else if (8'he5 == characterIndex) begin
            lengthsOut_229 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he6 == characterIndex) begin
              lengthsOut_230 <= _T_69;
            end
          end else if (8'he6 == characterIndex) begin
            lengthsOut_230 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he7 == characterIndex) begin
              lengthsOut_231 <= _T_69;
            end
          end else if (8'he7 == characterIndex) begin
            lengthsOut_231 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he8 == characterIndex) begin
              lengthsOut_232 <= _T_69;
            end
          end else if (8'he8 == characterIndex) begin
            lengthsOut_232 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'he9 == characterIndex) begin
              lengthsOut_233 <= _T_69;
            end
          end else if (8'he9 == characterIndex) begin
            lengthsOut_233 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hea == characterIndex) begin
              lengthsOut_234 <= _T_69;
            end
          end else if (8'hea == characterIndex) begin
            lengthsOut_234 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'heb == characterIndex) begin
              lengthsOut_235 <= _T_69;
            end
          end else if (8'heb == characterIndex) begin
            lengthsOut_235 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hec == characterIndex) begin
              lengthsOut_236 <= _T_69;
            end
          end else if (8'hec == characterIndex) begin
            lengthsOut_236 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hed == characterIndex) begin
              lengthsOut_237 <= _T_69;
            end
          end else if (8'hed == characterIndex) begin
            lengthsOut_237 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hee == characterIndex) begin
              lengthsOut_238 <= _T_69;
            end
          end else if (8'hee == characterIndex) begin
            lengthsOut_238 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hef == characterIndex) begin
              lengthsOut_239 <= _T_69;
            end
          end else if (8'hef == characterIndex) begin
            lengthsOut_239 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf0 == characterIndex) begin
              lengthsOut_240 <= _T_69;
            end
          end else if (8'hf0 == characterIndex) begin
            lengthsOut_240 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf1 == characterIndex) begin
              lengthsOut_241 <= _T_69;
            end
          end else if (8'hf1 == characterIndex) begin
            lengthsOut_241 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf2 == characterIndex) begin
              lengthsOut_242 <= _T_69;
            end
          end else if (8'hf2 == characterIndex) begin
            lengthsOut_242 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf3 == characterIndex) begin
              lengthsOut_243 <= _T_69;
            end
          end else if (8'hf3 == characterIndex) begin
            lengthsOut_243 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf4 == characterIndex) begin
              lengthsOut_244 <= _T_69;
            end
          end else if (8'hf4 == characterIndex) begin
            lengthsOut_244 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf5 == characterIndex) begin
              lengthsOut_245 <= _T_69;
            end
          end else if (8'hf5 == characterIndex) begin
            lengthsOut_245 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf6 == characterIndex) begin
              lengthsOut_246 <= _T_69;
            end
          end else if (8'hf6 == characterIndex) begin
            lengthsOut_246 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf7 == characterIndex) begin
              lengthsOut_247 <= _T_69;
            end
          end else if (8'hf7 == characterIndex) begin
            lengthsOut_247 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf8 == characterIndex) begin
              lengthsOut_248 <= _T_69;
            end
          end else if (8'hf8 == characterIndex) begin
            lengthsOut_248 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hf9 == characterIndex) begin
              lengthsOut_249 <= _T_69;
            end
          end else if (8'hf9 == characterIndex) begin
            lengthsOut_249 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hfa == characterIndex) begin
              lengthsOut_250 <= _T_69;
            end
          end else if (8'hfa == characterIndex) begin
            lengthsOut_250 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hfb == characterIndex) begin
              lengthsOut_251 <= _T_69;
            end
          end else if (8'hfb == characterIndex) begin
            lengthsOut_251 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hfc == characterIndex) begin
              lengthsOut_252 <= _T_69;
            end
          end else if (8'hfc == characterIndex) begin
            lengthsOut_252 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hfd == characterIndex) begin
              lengthsOut_253 <= _T_69;
            end
          end else if (8'hfd == characterIndex) begin
            lengthsOut_253 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hfe == characterIndex) begin
              lengthsOut_254 <= _T_69;
            end
          end else if (8'hfe == characterIndex) begin
            lengthsOut_254 <= _GEN_2550;
          end
        end
      end
    end
    if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (!(_T_30)) begin
          if (_T_66) begin
            if (8'hff == characterIndex) begin
              lengthsOut_255 <= _T_69;
            end
          end else if (8'hff == characterIndex) begin
            lengthsOut_255 <= _GEN_2550;
          end
        end
      end
    end
    if (reset) begin
      characterIndex <= 8'h0;
    end else if (_T_6) begin
      if (io_start) begin
        characterIndex <= 8'h0;
      end
    end else if (_T_9) begin
      if (_T_29) begin
        characterIndex <= 8'h0;
      end else begin
        characterIndex <= _T_12;
      end
    end else if (_T_30) begin
      if (_T_29) begin
        characterIndex <= 8'h0;
      end else if (!(_T_35)) begin
        characterIndex <= _T_12;
      end
    end else begin
      characterIndex <= _T_12;
    end
    if (reset) begin
      nodes <= 9'h0;
    end else if (_T_6) begin
      if (io_start) begin
        nodes <= io_inputs_validNodesOut;
      end
    end
    if (reset) begin
      characterDepth <= 4'h0;
    end else if (_T_6) begin
      if (io_start) begin
        characterDepth <= 4'h1;
      end
    end else if (!(_T_9)) begin
      if (_T_30) begin
        if (_T_35) begin
          if (5'h1f == characterIndex[4:0]) begin
            characterDepth <= depths_31;
          end else if (5'h1e == characterIndex[4:0]) begin
            characterDepth <= depths_30;
          end else if (5'h1d == characterIndex[4:0]) begin
            characterDepth <= depths_29;
          end else if (5'h1c == characterIndex[4:0]) begin
            characterDepth <= depths_28;
          end else if (5'h1b == characterIndex[4:0]) begin
            characterDepth <= depths_27;
          end else if (5'h1a == characterIndex[4:0]) begin
            characterDepth <= depths_26;
          end else if (5'h19 == characterIndex[4:0]) begin
            characterDepth <= depths_25;
          end else if (5'h18 == characterIndex[4:0]) begin
            characterDepth <= depths_24;
          end else if (5'h17 == characterIndex[4:0]) begin
            characterDepth <= depths_23;
          end else if (5'h16 == characterIndex[4:0]) begin
            characterDepth <= depths_22;
          end else if (5'h15 == characterIndex[4:0]) begin
            characterDepth <= depths_21;
          end else if (5'h14 == characterIndex[4:0]) begin
            characterDepth <= depths_20;
          end else if (5'h13 == characterIndex[4:0]) begin
            characterDepth <= depths_19;
          end else if (5'h12 == characterIndex[4:0]) begin
            characterDepth <= depths_18;
          end else if (5'h11 == characterIndex[4:0]) begin
            characterDepth <= depths_17;
          end else if (5'h10 == characterIndex[4:0]) begin
            characterDepth <= depths_16;
          end else if (5'hf == characterIndex[4:0]) begin
            characterDepth <= depths_15;
          end else if (5'he == characterIndex[4:0]) begin
            characterDepth <= depths_14;
          end else if (5'hd == characterIndex[4:0]) begin
            characterDepth <= depths_13;
          end else if (5'hc == characterIndex[4:0]) begin
            characterDepth <= depths_12;
          end else if (5'hb == characterIndex[4:0]) begin
            characterDepth <= depths_11;
          end else if (5'ha == characterIndex[4:0]) begin
            characterDepth <= depths_10;
          end else if (5'h9 == characterIndex[4:0]) begin
            characterDepth <= depths_9;
          end else if (5'h8 == characterIndex[4:0]) begin
            characterDepth <= depths_8;
          end else if (5'h7 == characterIndex[4:0]) begin
            characterDepth <= depths_7;
          end else if (5'h6 == characterIndex[4:0]) begin
            characterDepth <= depths_6;
          end else if (5'h5 == characterIndex[4:0]) begin
            characterDepth <= depths_5;
          end else if (5'h4 == characterIndex[4:0]) begin
            characterDepth <= depths_4;
          end else if (5'h3 == characterIndex[4:0]) begin
            characterDepth <= depths_3;
          end else if (5'h2 == characterIndex[4:0]) begin
            characterDepth <= depths_2;
          end else if (5'h1 == characterIndex[4:0]) begin
            characterDepth <= depths_1;
          end else begin
            characterDepth <= depths_0;
          end
        end
      end
    end
    if (reset) begin
      codeword <= 16'h0;
    end else begin
      codeword <= _GEN_7835[15:0];
    end
    if (reset) begin
      escapeCodeword <= 16'h0;
    end else if (!(_T_6)) begin
      if (!(_T_9)) begin
        if (_T_30) begin
          if (!(_T_35)) begin
            if (_GEN_182[8]) begin
              escapeCodeword <= codeword;
            end
          end
        end
      end
    end
    if (reset) begin
      escapeCharacterLength <= 4'h0;
    end else if (_T_6) begin
      if (io_start) begin
        escapeCharacterLength <= 4'h0;
      end
    end else if (!(_T_9)) begin
      if (_T_30) begin
        if (!(_T_35)) begin
          if (_GEN_182[8]) begin
            escapeCharacterLength <= characterDepth;
          end
        end
      end
    end
  end
endmodule
module compressorOutput(
  input         clock,
  input         reset,
  input         io_start,
  output [11:0] io_dataIn_0_currentByteOut,
  input  [7:0]  io_dataIn_0_dataIn_0,
  input         io_dataIn_0_valid,
  output        io_dataIn_0_ready,
  input  [23:0] io_inputs_codewords_0,
  input  [23:0] io_inputs_codewords_1,
  input  [23:0] io_inputs_codewords_2,
  input  [23:0] io_inputs_codewords_3,
  input  [23:0] io_inputs_codewords_4,
  input  [23:0] io_inputs_codewords_5,
  input  [23:0] io_inputs_codewords_6,
  input  [23:0] io_inputs_codewords_7,
  input  [23:0] io_inputs_codewords_8,
  input  [23:0] io_inputs_codewords_9,
  input  [23:0] io_inputs_codewords_10,
  input  [23:0] io_inputs_codewords_11,
  input  [23:0] io_inputs_codewords_12,
  input  [23:0] io_inputs_codewords_13,
  input  [23:0] io_inputs_codewords_14,
  input  [23:0] io_inputs_codewords_15,
  input  [23:0] io_inputs_codewords_16,
  input  [23:0] io_inputs_codewords_17,
  input  [23:0] io_inputs_codewords_18,
  input  [23:0] io_inputs_codewords_19,
  input  [23:0] io_inputs_codewords_20,
  input  [23:0] io_inputs_codewords_21,
  input  [23:0] io_inputs_codewords_22,
  input  [23:0] io_inputs_codewords_23,
  input  [23:0] io_inputs_codewords_24,
  input  [23:0] io_inputs_codewords_25,
  input  [23:0] io_inputs_codewords_26,
  input  [23:0] io_inputs_codewords_27,
  input  [23:0] io_inputs_codewords_28,
  input  [23:0] io_inputs_codewords_29,
  input  [23:0] io_inputs_codewords_30,
  input  [23:0] io_inputs_codewords_31,
  input  [23:0] io_inputs_codewords_32,
  input  [23:0] io_inputs_codewords_33,
  input  [23:0] io_inputs_codewords_34,
  input  [23:0] io_inputs_codewords_35,
  input  [23:0] io_inputs_codewords_36,
  input  [23:0] io_inputs_codewords_37,
  input  [23:0] io_inputs_codewords_38,
  input  [23:0] io_inputs_codewords_39,
  input  [23:0] io_inputs_codewords_40,
  input  [23:0] io_inputs_codewords_41,
  input  [23:0] io_inputs_codewords_42,
  input  [23:0] io_inputs_codewords_43,
  input  [23:0] io_inputs_codewords_44,
  input  [23:0] io_inputs_codewords_45,
  input  [23:0] io_inputs_codewords_46,
  input  [23:0] io_inputs_codewords_47,
  input  [23:0] io_inputs_codewords_48,
  input  [23:0] io_inputs_codewords_49,
  input  [23:0] io_inputs_codewords_50,
  input  [23:0] io_inputs_codewords_51,
  input  [23:0] io_inputs_codewords_52,
  input  [23:0] io_inputs_codewords_53,
  input  [23:0] io_inputs_codewords_54,
  input  [23:0] io_inputs_codewords_55,
  input  [23:0] io_inputs_codewords_56,
  input  [23:0] io_inputs_codewords_57,
  input  [23:0] io_inputs_codewords_58,
  input  [23:0] io_inputs_codewords_59,
  input  [23:0] io_inputs_codewords_60,
  input  [23:0] io_inputs_codewords_61,
  input  [23:0] io_inputs_codewords_62,
  input  [23:0] io_inputs_codewords_63,
  input  [23:0] io_inputs_codewords_64,
  input  [23:0] io_inputs_codewords_65,
  input  [23:0] io_inputs_codewords_66,
  input  [23:0] io_inputs_codewords_67,
  input  [23:0] io_inputs_codewords_68,
  input  [23:0] io_inputs_codewords_69,
  input  [23:0] io_inputs_codewords_70,
  input  [23:0] io_inputs_codewords_71,
  input  [23:0] io_inputs_codewords_72,
  input  [23:0] io_inputs_codewords_73,
  input  [23:0] io_inputs_codewords_74,
  input  [23:0] io_inputs_codewords_75,
  input  [23:0] io_inputs_codewords_76,
  input  [23:0] io_inputs_codewords_77,
  input  [23:0] io_inputs_codewords_78,
  input  [23:0] io_inputs_codewords_79,
  input  [23:0] io_inputs_codewords_80,
  input  [23:0] io_inputs_codewords_81,
  input  [23:0] io_inputs_codewords_82,
  input  [23:0] io_inputs_codewords_83,
  input  [23:0] io_inputs_codewords_84,
  input  [23:0] io_inputs_codewords_85,
  input  [23:0] io_inputs_codewords_86,
  input  [23:0] io_inputs_codewords_87,
  input  [23:0] io_inputs_codewords_88,
  input  [23:0] io_inputs_codewords_89,
  input  [23:0] io_inputs_codewords_90,
  input  [23:0] io_inputs_codewords_91,
  input  [23:0] io_inputs_codewords_92,
  input  [23:0] io_inputs_codewords_93,
  input  [23:0] io_inputs_codewords_94,
  input  [23:0] io_inputs_codewords_95,
  input  [23:0] io_inputs_codewords_96,
  input  [23:0] io_inputs_codewords_97,
  input  [23:0] io_inputs_codewords_98,
  input  [23:0] io_inputs_codewords_99,
  input  [23:0] io_inputs_codewords_100,
  input  [23:0] io_inputs_codewords_101,
  input  [23:0] io_inputs_codewords_102,
  input  [23:0] io_inputs_codewords_103,
  input  [23:0] io_inputs_codewords_104,
  input  [23:0] io_inputs_codewords_105,
  input  [23:0] io_inputs_codewords_106,
  input  [23:0] io_inputs_codewords_107,
  input  [23:0] io_inputs_codewords_108,
  input  [23:0] io_inputs_codewords_109,
  input  [23:0] io_inputs_codewords_110,
  input  [23:0] io_inputs_codewords_111,
  input  [23:0] io_inputs_codewords_112,
  input  [23:0] io_inputs_codewords_113,
  input  [23:0] io_inputs_codewords_114,
  input  [23:0] io_inputs_codewords_115,
  input  [23:0] io_inputs_codewords_116,
  input  [23:0] io_inputs_codewords_117,
  input  [23:0] io_inputs_codewords_118,
  input  [23:0] io_inputs_codewords_119,
  input  [23:0] io_inputs_codewords_120,
  input  [23:0] io_inputs_codewords_121,
  input  [23:0] io_inputs_codewords_122,
  input  [23:0] io_inputs_codewords_123,
  input  [23:0] io_inputs_codewords_124,
  input  [23:0] io_inputs_codewords_125,
  input  [23:0] io_inputs_codewords_126,
  input  [23:0] io_inputs_codewords_127,
  input  [23:0] io_inputs_codewords_128,
  input  [23:0] io_inputs_codewords_129,
  input  [23:0] io_inputs_codewords_130,
  input  [23:0] io_inputs_codewords_131,
  input  [23:0] io_inputs_codewords_132,
  input  [23:0] io_inputs_codewords_133,
  input  [23:0] io_inputs_codewords_134,
  input  [23:0] io_inputs_codewords_135,
  input  [23:0] io_inputs_codewords_136,
  input  [23:0] io_inputs_codewords_137,
  input  [23:0] io_inputs_codewords_138,
  input  [23:0] io_inputs_codewords_139,
  input  [23:0] io_inputs_codewords_140,
  input  [23:0] io_inputs_codewords_141,
  input  [23:0] io_inputs_codewords_142,
  input  [23:0] io_inputs_codewords_143,
  input  [23:0] io_inputs_codewords_144,
  input  [23:0] io_inputs_codewords_145,
  input  [23:0] io_inputs_codewords_146,
  input  [23:0] io_inputs_codewords_147,
  input  [23:0] io_inputs_codewords_148,
  input  [23:0] io_inputs_codewords_149,
  input  [23:0] io_inputs_codewords_150,
  input  [23:0] io_inputs_codewords_151,
  input  [23:0] io_inputs_codewords_152,
  input  [23:0] io_inputs_codewords_153,
  input  [23:0] io_inputs_codewords_154,
  input  [23:0] io_inputs_codewords_155,
  input  [23:0] io_inputs_codewords_156,
  input  [23:0] io_inputs_codewords_157,
  input  [23:0] io_inputs_codewords_158,
  input  [23:0] io_inputs_codewords_159,
  input  [23:0] io_inputs_codewords_160,
  input  [23:0] io_inputs_codewords_161,
  input  [23:0] io_inputs_codewords_162,
  input  [23:0] io_inputs_codewords_163,
  input  [23:0] io_inputs_codewords_164,
  input  [23:0] io_inputs_codewords_165,
  input  [23:0] io_inputs_codewords_166,
  input  [23:0] io_inputs_codewords_167,
  input  [23:0] io_inputs_codewords_168,
  input  [23:0] io_inputs_codewords_169,
  input  [23:0] io_inputs_codewords_170,
  input  [23:0] io_inputs_codewords_171,
  input  [23:0] io_inputs_codewords_172,
  input  [23:0] io_inputs_codewords_173,
  input  [23:0] io_inputs_codewords_174,
  input  [23:0] io_inputs_codewords_175,
  input  [23:0] io_inputs_codewords_176,
  input  [23:0] io_inputs_codewords_177,
  input  [23:0] io_inputs_codewords_178,
  input  [23:0] io_inputs_codewords_179,
  input  [23:0] io_inputs_codewords_180,
  input  [23:0] io_inputs_codewords_181,
  input  [23:0] io_inputs_codewords_182,
  input  [23:0] io_inputs_codewords_183,
  input  [23:0] io_inputs_codewords_184,
  input  [23:0] io_inputs_codewords_185,
  input  [23:0] io_inputs_codewords_186,
  input  [23:0] io_inputs_codewords_187,
  input  [23:0] io_inputs_codewords_188,
  input  [23:0] io_inputs_codewords_189,
  input  [23:0] io_inputs_codewords_190,
  input  [23:0] io_inputs_codewords_191,
  input  [23:0] io_inputs_codewords_192,
  input  [23:0] io_inputs_codewords_193,
  input  [23:0] io_inputs_codewords_194,
  input  [23:0] io_inputs_codewords_195,
  input  [23:0] io_inputs_codewords_196,
  input  [23:0] io_inputs_codewords_197,
  input  [23:0] io_inputs_codewords_198,
  input  [23:0] io_inputs_codewords_199,
  input  [23:0] io_inputs_codewords_200,
  input  [23:0] io_inputs_codewords_201,
  input  [23:0] io_inputs_codewords_202,
  input  [23:0] io_inputs_codewords_203,
  input  [23:0] io_inputs_codewords_204,
  input  [23:0] io_inputs_codewords_205,
  input  [23:0] io_inputs_codewords_206,
  input  [23:0] io_inputs_codewords_207,
  input  [23:0] io_inputs_codewords_208,
  input  [23:0] io_inputs_codewords_209,
  input  [23:0] io_inputs_codewords_210,
  input  [23:0] io_inputs_codewords_211,
  input  [23:0] io_inputs_codewords_212,
  input  [23:0] io_inputs_codewords_213,
  input  [23:0] io_inputs_codewords_214,
  input  [23:0] io_inputs_codewords_215,
  input  [23:0] io_inputs_codewords_216,
  input  [23:0] io_inputs_codewords_217,
  input  [23:0] io_inputs_codewords_218,
  input  [23:0] io_inputs_codewords_219,
  input  [23:0] io_inputs_codewords_220,
  input  [23:0] io_inputs_codewords_221,
  input  [23:0] io_inputs_codewords_222,
  input  [23:0] io_inputs_codewords_223,
  input  [23:0] io_inputs_codewords_224,
  input  [23:0] io_inputs_codewords_225,
  input  [23:0] io_inputs_codewords_226,
  input  [23:0] io_inputs_codewords_227,
  input  [23:0] io_inputs_codewords_228,
  input  [23:0] io_inputs_codewords_229,
  input  [23:0] io_inputs_codewords_230,
  input  [23:0] io_inputs_codewords_231,
  input  [23:0] io_inputs_codewords_232,
  input  [23:0] io_inputs_codewords_233,
  input  [23:0] io_inputs_codewords_234,
  input  [23:0] io_inputs_codewords_235,
  input  [23:0] io_inputs_codewords_236,
  input  [23:0] io_inputs_codewords_237,
  input  [23:0] io_inputs_codewords_238,
  input  [23:0] io_inputs_codewords_239,
  input  [23:0] io_inputs_codewords_240,
  input  [23:0] io_inputs_codewords_241,
  input  [23:0] io_inputs_codewords_242,
  input  [23:0] io_inputs_codewords_243,
  input  [23:0] io_inputs_codewords_244,
  input  [23:0] io_inputs_codewords_245,
  input  [23:0] io_inputs_codewords_246,
  input  [23:0] io_inputs_codewords_247,
  input  [23:0] io_inputs_codewords_248,
  input  [23:0] io_inputs_codewords_249,
  input  [23:0] io_inputs_codewords_250,
  input  [23:0] io_inputs_codewords_251,
  input  [23:0] io_inputs_codewords_252,
  input  [23:0] io_inputs_codewords_253,
  input  [23:0] io_inputs_codewords_254,
  input  [23:0] io_inputs_codewords_255,
  input  [4:0]  io_inputs_lengths_0,
  input  [4:0]  io_inputs_lengths_1,
  input  [4:0]  io_inputs_lengths_2,
  input  [4:0]  io_inputs_lengths_3,
  input  [4:0]  io_inputs_lengths_4,
  input  [4:0]  io_inputs_lengths_5,
  input  [4:0]  io_inputs_lengths_6,
  input  [4:0]  io_inputs_lengths_7,
  input  [4:0]  io_inputs_lengths_8,
  input  [4:0]  io_inputs_lengths_9,
  input  [4:0]  io_inputs_lengths_10,
  input  [4:0]  io_inputs_lengths_11,
  input  [4:0]  io_inputs_lengths_12,
  input  [4:0]  io_inputs_lengths_13,
  input  [4:0]  io_inputs_lengths_14,
  input  [4:0]  io_inputs_lengths_15,
  input  [4:0]  io_inputs_lengths_16,
  input  [4:0]  io_inputs_lengths_17,
  input  [4:0]  io_inputs_lengths_18,
  input  [4:0]  io_inputs_lengths_19,
  input  [4:0]  io_inputs_lengths_20,
  input  [4:0]  io_inputs_lengths_21,
  input  [4:0]  io_inputs_lengths_22,
  input  [4:0]  io_inputs_lengths_23,
  input  [4:0]  io_inputs_lengths_24,
  input  [4:0]  io_inputs_lengths_25,
  input  [4:0]  io_inputs_lengths_26,
  input  [4:0]  io_inputs_lengths_27,
  input  [4:0]  io_inputs_lengths_28,
  input  [4:0]  io_inputs_lengths_29,
  input  [4:0]  io_inputs_lengths_30,
  input  [4:0]  io_inputs_lengths_31,
  input  [4:0]  io_inputs_lengths_32,
  input  [4:0]  io_inputs_lengths_33,
  input  [4:0]  io_inputs_lengths_34,
  input  [4:0]  io_inputs_lengths_35,
  input  [4:0]  io_inputs_lengths_36,
  input  [4:0]  io_inputs_lengths_37,
  input  [4:0]  io_inputs_lengths_38,
  input  [4:0]  io_inputs_lengths_39,
  input  [4:0]  io_inputs_lengths_40,
  input  [4:0]  io_inputs_lengths_41,
  input  [4:0]  io_inputs_lengths_42,
  input  [4:0]  io_inputs_lengths_43,
  input  [4:0]  io_inputs_lengths_44,
  input  [4:0]  io_inputs_lengths_45,
  input  [4:0]  io_inputs_lengths_46,
  input  [4:0]  io_inputs_lengths_47,
  input  [4:0]  io_inputs_lengths_48,
  input  [4:0]  io_inputs_lengths_49,
  input  [4:0]  io_inputs_lengths_50,
  input  [4:0]  io_inputs_lengths_51,
  input  [4:0]  io_inputs_lengths_52,
  input  [4:0]  io_inputs_lengths_53,
  input  [4:0]  io_inputs_lengths_54,
  input  [4:0]  io_inputs_lengths_55,
  input  [4:0]  io_inputs_lengths_56,
  input  [4:0]  io_inputs_lengths_57,
  input  [4:0]  io_inputs_lengths_58,
  input  [4:0]  io_inputs_lengths_59,
  input  [4:0]  io_inputs_lengths_60,
  input  [4:0]  io_inputs_lengths_61,
  input  [4:0]  io_inputs_lengths_62,
  input  [4:0]  io_inputs_lengths_63,
  input  [4:0]  io_inputs_lengths_64,
  input  [4:0]  io_inputs_lengths_65,
  input  [4:0]  io_inputs_lengths_66,
  input  [4:0]  io_inputs_lengths_67,
  input  [4:0]  io_inputs_lengths_68,
  input  [4:0]  io_inputs_lengths_69,
  input  [4:0]  io_inputs_lengths_70,
  input  [4:0]  io_inputs_lengths_71,
  input  [4:0]  io_inputs_lengths_72,
  input  [4:0]  io_inputs_lengths_73,
  input  [4:0]  io_inputs_lengths_74,
  input  [4:0]  io_inputs_lengths_75,
  input  [4:0]  io_inputs_lengths_76,
  input  [4:0]  io_inputs_lengths_77,
  input  [4:0]  io_inputs_lengths_78,
  input  [4:0]  io_inputs_lengths_79,
  input  [4:0]  io_inputs_lengths_80,
  input  [4:0]  io_inputs_lengths_81,
  input  [4:0]  io_inputs_lengths_82,
  input  [4:0]  io_inputs_lengths_83,
  input  [4:0]  io_inputs_lengths_84,
  input  [4:0]  io_inputs_lengths_85,
  input  [4:0]  io_inputs_lengths_86,
  input  [4:0]  io_inputs_lengths_87,
  input  [4:0]  io_inputs_lengths_88,
  input  [4:0]  io_inputs_lengths_89,
  input  [4:0]  io_inputs_lengths_90,
  input  [4:0]  io_inputs_lengths_91,
  input  [4:0]  io_inputs_lengths_92,
  input  [4:0]  io_inputs_lengths_93,
  input  [4:0]  io_inputs_lengths_94,
  input  [4:0]  io_inputs_lengths_95,
  input  [4:0]  io_inputs_lengths_96,
  input  [4:0]  io_inputs_lengths_97,
  input  [4:0]  io_inputs_lengths_98,
  input  [4:0]  io_inputs_lengths_99,
  input  [4:0]  io_inputs_lengths_100,
  input  [4:0]  io_inputs_lengths_101,
  input  [4:0]  io_inputs_lengths_102,
  input  [4:0]  io_inputs_lengths_103,
  input  [4:0]  io_inputs_lengths_104,
  input  [4:0]  io_inputs_lengths_105,
  input  [4:0]  io_inputs_lengths_106,
  input  [4:0]  io_inputs_lengths_107,
  input  [4:0]  io_inputs_lengths_108,
  input  [4:0]  io_inputs_lengths_109,
  input  [4:0]  io_inputs_lengths_110,
  input  [4:0]  io_inputs_lengths_111,
  input  [4:0]  io_inputs_lengths_112,
  input  [4:0]  io_inputs_lengths_113,
  input  [4:0]  io_inputs_lengths_114,
  input  [4:0]  io_inputs_lengths_115,
  input  [4:0]  io_inputs_lengths_116,
  input  [4:0]  io_inputs_lengths_117,
  input  [4:0]  io_inputs_lengths_118,
  input  [4:0]  io_inputs_lengths_119,
  input  [4:0]  io_inputs_lengths_120,
  input  [4:0]  io_inputs_lengths_121,
  input  [4:0]  io_inputs_lengths_122,
  input  [4:0]  io_inputs_lengths_123,
  input  [4:0]  io_inputs_lengths_124,
  input  [4:0]  io_inputs_lengths_125,
  input  [4:0]  io_inputs_lengths_126,
  input  [4:0]  io_inputs_lengths_127,
  input  [4:0]  io_inputs_lengths_128,
  input  [4:0]  io_inputs_lengths_129,
  input  [4:0]  io_inputs_lengths_130,
  input  [4:0]  io_inputs_lengths_131,
  input  [4:0]  io_inputs_lengths_132,
  input  [4:0]  io_inputs_lengths_133,
  input  [4:0]  io_inputs_lengths_134,
  input  [4:0]  io_inputs_lengths_135,
  input  [4:0]  io_inputs_lengths_136,
  input  [4:0]  io_inputs_lengths_137,
  input  [4:0]  io_inputs_lengths_138,
  input  [4:0]  io_inputs_lengths_139,
  input  [4:0]  io_inputs_lengths_140,
  input  [4:0]  io_inputs_lengths_141,
  input  [4:0]  io_inputs_lengths_142,
  input  [4:0]  io_inputs_lengths_143,
  input  [4:0]  io_inputs_lengths_144,
  input  [4:0]  io_inputs_lengths_145,
  input  [4:0]  io_inputs_lengths_146,
  input  [4:0]  io_inputs_lengths_147,
  input  [4:0]  io_inputs_lengths_148,
  input  [4:0]  io_inputs_lengths_149,
  input  [4:0]  io_inputs_lengths_150,
  input  [4:0]  io_inputs_lengths_151,
  input  [4:0]  io_inputs_lengths_152,
  input  [4:0]  io_inputs_lengths_153,
  input  [4:0]  io_inputs_lengths_154,
  input  [4:0]  io_inputs_lengths_155,
  input  [4:0]  io_inputs_lengths_156,
  input  [4:0]  io_inputs_lengths_157,
  input  [4:0]  io_inputs_lengths_158,
  input  [4:0]  io_inputs_lengths_159,
  input  [4:0]  io_inputs_lengths_160,
  input  [4:0]  io_inputs_lengths_161,
  input  [4:0]  io_inputs_lengths_162,
  input  [4:0]  io_inputs_lengths_163,
  input  [4:0]  io_inputs_lengths_164,
  input  [4:0]  io_inputs_lengths_165,
  input  [4:0]  io_inputs_lengths_166,
  input  [4:0]  io_inputs_lengths_167,
  input  [4:0]  io_inputs_lengths_168,
  input  [4:0]  io_inputs_lengths_169,
  input  [4:0]  io_inputs_lengths_170,
  input  [4:0]  io_inputs_lengths_171,
  input  [4:0]  io_inputs_lengths_172,
  input  [4:0]  io_inputs_lengths_173,
  input  [4:0]  io_inputs_lengths_174,
  input  [4:0]  io_inputs_lengths_175,
  input  [4:0]  io_inputs_lengths_176,
  input  [4:0]  io_inputs_lengths_177,
  input  [4:0]  io_inputs_lengths_178,
  input  [4:0]  io_inputs_lengths_179,
  input  [4:0]  io_inputs_lengths_180,
  input  [4:0]  io_inputs_lengths_181,
  input  [4:0]  io_inputs_lengths_182,
  input  [4:0]  io_inputs_lengths_183,
  input  [4:0]  io_inputs_lengths_184,
  input  [4:0]  io_inputs_lengths_185,
  input  [4:0]  io_inputs_lengths_186,
  input  [4:0]  io_inputs_lengths_187,
  input  [4:0]  io_inputs_lengths_188,
  input  [4:0]  io_inputs_lengths_189,
  input  [4:0]  io_inputs_lengths_190,
  input  [4:0]  io_inputs_lengths_191,
  input  [4:0]  io_inputs_lengths_192,
  input  [4:0]  io_inputs_lengths_193,
  input  [4:0]  io_inputs_lengths_194,
  input  [4:0]  io_inputs_lengths_195,
  input  [4:0]  io_inputs_lengths_196,
  input  [4:0]  io_inputs_lengths_197,
  input  [4:0]  io_inputs_lengths_198,
  input  [4:0]  io_inputs_lengths_199,
  input  [4:0]  io_inputs_lengths_200,
  input  [4:0]  io_inputs_lengths_201,
  input  [4:0]  io_inputs_lengths_202,
  input  [4:0]  io_inputs_lengths_203,
  input  [4:0]  io_inputs_lengths_204,
  input  [4:0]  io_inputs_lengths_205,
  input  [4:0]  io_inputs_lengths_206,
  input  [4:0]  io_inputs_lengths_207,
  input  [4:0]  io_inputs_lengths_208,
  input  [4:0]  io_inputs_lengths_209,
  input  [4:0]  io_inputs_lengths_210,
  input  [4:0]  io_inputs_lengths_211,
  input  [4:0]  io_inputs_lengths_212,
  input  [4:0]  io_inputs_lengths_213,
  input  [4:0]  io_inputs_lengths_214,
  input  [4:0]  io_inputs_lengths_215,
  input  [4:0]  io_inputs_lengths_216,
  input  [4:0]  io_inputs_lengths_217,
  input  [4:0]  io_inputs_lengths_218,
  input  [4:0]  io_inputs_lengths_219,
  input  [4:0]  io_inputs_lengths_220,
  input  [4:0]  io_inputs_lengths_221,
  input  [4:0]  io_inputs_lengths_222,
  input  [4:0]  io_inputs_lengths_223,
  input  [4:0]  io_inputs_lengths_224,
  input  [4:0]  io_inputs_lengths_225,
  input  [4:0]  io_inputs_lengths_226,
  input  [4:0]  io_inputs_lengths_227,
  input  [4:0]  io_inputs_lengths_228,
  input  [4:0]  io_inputs_lengths_229,
  input  [4:0]  io_inputs_lengths_230,
  input  [4:0]  io_inputs_lengths_231,
  input  [4:0]  io_inputs_lengths_232,
  input  [4:0]  io_inputs_lengths_233,
  input  [4:0]  io_inputs_lengths_234,
  input  [4:0]  io_inputs_lengths_235,
  input  [4:0]  io_inputs_lengths_236,
  input  [4:0]  io_inputs_lengths_237,
  input  [4:0]  io_inputs_lengths_238,
  input  [4:0]  io_inputs_lengths_239,
  input  [4:0]  io_inputs_lengths_240,
  input  [4:0]  io_inputs_lengths_241,
  input  [4:0]  io_inputs_lengths_242,
  input  [4:0]  io_inputs_lengths_243,
  input  [4:0]  io_inputs_lengths_244,
  input  [4:0]  io_inputs_lengths_245,
  input  [4:0]  io_inputs_lengths_246,
  input  [4:0]  io_inputs_lengths_247,
  input  [4:0]  io_inputs_lengths_248,
  input  [4:0]  io_inputs_lengths_249,
  input  [4:0]  io_inputs_lengths_250,
  input  [4:0]  io_inputs_lengths_251,
  input  [4:0]  io_inputs_lengths_252,
  input  [4:0]  io_inputs_lengths_253,
  input  [4:0]  io_inputs_lengths_254,
  input  [4:0]  io_inputs_lengths_255,
  input  [8:0]  io_inputs_charactersOut_0,
  input  [8:0]  io_inputs_charactersOut_1,
  input  [8:0]  io_inputs_charactersOut_2,
  input  [8:0]  io_inputs_charactersOut_3,
  input  [8:0]  io_inputs_charactersOut_4,
  input  [8:0]  io_inputs_charactersOut_5,
  input  [8:0]  io_inputs_charactersOut_6,
  input  [8:0]  io_inputs_charactersOut_7,
  input  [8:0]  io_inputs_charactersOut_8,
  input  [8:0]  io_inputs_charactersOut_9,
  input  [8:0]  io_inputs_charactersOut_10,
  input  [8:0]  io_inputs_charactersOut_11,
  input  [8:0]  io_inputs_charactersOut_12,
  input  [8:0]  io_inputs_charactersOut_13,
  input  [8:0]  io_inputs_charactersOut_14,
  input  [8:0]  io_inputs_charactersOut_15,
  input  [8:0]  io_inputs_charactersOut_16,
  input  [8:0]  io_inputs_charactersOut_17,
  input  [8:0]  io_inputs_charactersOut_18,
  input  [8:0]  io_inputs_charactersOut_19,
  input  [8:0]  io_inputs_charactersOut_20,
  input  [8:0]  io_inputs_charactersOut_21,
  input  [8:0]  io_inputs_charactersOut_22,
  input  [8:0]  io_inputs_charactersOut_23,
  input  [8:0]  io_inputs_charactersOut_24,
  input  [8:0]  io_inputs_charactersOut_25,
  input  [8:0]  io_inputs_charactersOut_26,
  input  [8:0]  io_inputs_charactersOut_27,
  input  [8:0]  io_inputs_charactersOut_28,
  input  [8:0]  io_inputs_charactersOut_29,
  input  [8:0]  io_inputs_charactersOut_30,
  input  [8:0]  io_inputs_charactersOut_31,
  input  [8:0]  io_inputs_nodes,
  input  [3:0]  io_inputs_escapeCharacterLength,
  input  [15:0] io_inputs_escapeCodeword,
  output [27:0] io_outputs_0_dataOut,
  output [4:0]  io_outputs_0_dataLength,
  output        io_outputs_0_valid,
  input         io_outputs_0_ready,
  output        io_finished
);
  wire [11:0] input_0_io_input_currentByteOut; // @[compressorOutput.scala 34:51]
  wire [7:0] input_0_io_input_dataIn_0; // @[compressorOutput.scala 34:51]
  wire  input_0_io_input_valid; // @[compressorOutput.scala 34:51]
  wire  input_0_io_input_ready; // @[compressorOutput.scala 34:51]
  wire [11:0] input_0_io_currentByte; // @[compressorOutput.scala 34:51]
  wire  input_0_io_dataOut_ready; // @[compressorOutput.scala 34:51]
  wire  input_0_io_dataOut_valid; // @[compressorOutput.scala 34:51]
  wire [7:0] input_0_io_dataOut_bits_0; // @[compressorOutput.scala 34:51]
  reg [1:0] state; // @[compressorOutput.scala 39:22]
  reg [31:0] _RAND_0;
  reg [12:0] iterations_0; // @[compressorOutput.scala 41:23]
  reg [31:0] _RAND_1;
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire [12:0] _GEN_1222 = {{4'd0}, io_inputs_nodes}; // @[compressorOutput.scala 87:26]
  wire  _T_2 = iterations_0 < _GEN_1222; // @[compressorOutput.scala 87:26]
  wire [8:0] _GEN_2 = 5'h1 == iterations_0[4:0] ? io_inputs_charactersOut_1 : io_inputs_charactersOut_0; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_3 = 5'h2 == iterations_0[4:0] ? io_inputs_charactersOut_2 : _GEN_2; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_4 = 5'h3 == iterations_0[4:0] ? io_inputs_charactersOut_3 : _GEN_3; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_5 = 5'h4 == iterations_0[4:0] ? io_inputs_charactersOut_4 : _GEN_4; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_6 = 5'h5 == iterations_0[4:0] ? io_inputs_charactersOut_5 : _GEN_5; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_7 = 5'h6 == iterations_0[4:0] ? io_inputs_charactersOut_6 : _GEN_6; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_8 = 5'h7 == iterations_0[4:0] ? io_inputs_charactersOut_7 : _GEN_7; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_9 = 5'h8 == iterations_0[4:0] ? io_inputs_charactersOut_8 : _GEN_8; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_10 = 5'h9 == iterations_0[4:0] ? io_inputs_charactersOut_9 : _GEN_9; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_11 = 5'ha == iterations_0[4:0] ? io_inputs_charactersOut_10 : _GEN_10; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_12 = 5'hb == iterations_0[4:0] ? io_inputs_charactersOut_11 : _GEN_11; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_13 = 5'hc == iterations_0[4:0] ? io_inputs_charactersOut_12 : _GEN_12; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_14 = 5'hd == iterations_0[4:0] ? io_inputs_charactersOut_13 : _GEN_13; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_15 = 5'he == iterations_0[4:0] ? io_inputs_charactersOut_14 : _GEN_14; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_16 = 5'hf == iterations_0[4:0] ? io_inputs_charactersOut_15 : _GEN_15; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_17 = 5'h10 == iterations_0[4:0] ? io_inputs_charactersOut_16 : _GEN_16; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_18 = 5'h11 == iterations_0[4:0] ? io_inputs_charactersOut_17 : _GEN_17; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_19 = 5'h12 == iterations_0[4:0] ? io_inputs_charactersOut_18 : _GEN_18; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_20 = 5'h13 == iterations_0[4:0] ? io_inputs_charactersOut_19 : _GEN_19; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_21 = 5'h14 == iterations_0[4:0] ? io_inputs_charactersOut_20 : _GEN_20; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_22 = 5'h15 == iterations_0[4:0] ? io_inputs_charactersOut_21 : _GEN_21; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_23 = 5'h16 == iterations_0[4:0] ? io_inputs_charactersOut_22 : _GEN_22; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_24 = 5'h17 == iterations_0[4:0] ? io_inputs_charactersOut_23 : _GEN_23; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_25 = 5'h18 == iterations_0[4:0] ? io_inputs_charactersOut_24 : _GEN_24; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_26 = 5'h19 == iterations_0[4:0] ? io_inputs_charactersOut_25 : _GEN_25; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_27 = 5'h1a == iterations_0[4:0] ? io_inputs_charactersOut_26 : _GEN_26; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_28 = 5'h1b == iterations_0[4:0] ? io_inputs_charactersOut_27 : _GEN_27; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_29 = 5'h1c == iterations_0[4:0] ? io_inputs_charactersOut_28 : _GEN_28; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_30 = 5'h1d == iterations_0[4:0] ? io_inputs_charactersOut_29 : _GEN_29; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_31 = 5'h1e == iterations_0[4:0] ? io_inputs_charactersOut_30 : _GEN_30; // @[compressorOutput.scala 89:49]
  wire [8:0] _GEN_32 = 5'h1f == iterations_0[4:0] ? io_inputs_charactersOut_31 : _GEN_31; // @[compressorOutput.scala 89:49]
  wire [27:0] _T_9 = {_GEN_32,io_inputs_escapeCodeword[14:0],io_inputs_escapeCharacterLength}; // @[Cat.scala 29:58]
  wire [23:0] _GEN_98 = 8'h1 == _GEN_32[7:0] ? io_inputs_codewords_1 : io_inputs_codewords_0; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_99 = 8'h2 == _GEN_32[7:0] ? io_inputs_codewords_2 : _GEN_98; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_100 = 8'h3 == _GEN_32[7:0] ? io_inputs_codewords_3 : _GEN_99; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_101 = 8'h4 == _GEN_32[7:0] ? io_inputs_codewords_4 : _GEN_100; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_102 = 8'h5 == _GEN_32[7:0] ? io_inputs_codewords_5 : _GEN_101; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_103 = 8'h6 == _GEN_32[7:0] ? io_inputs_codewords_6 : _GEN_102; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_104 = 8'h7 == _GEN_32[7:0] ? io_inputs_codewords_7 : _GEN_103; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_105 = 8'h8 == _GEN_32[7:0] ? io_inputs_codewords_8 : _GEN_104; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_106 = 8'h9 == _GEN_32[7:0] ? io_inputs_codewords_9 : _GEN_105; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_107 = 8'ha == _GEN_32[7:0] ? io_inputs_codewords_10 : _GEN_106; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_108 = 8'hb == _GEN_32[7:0] ? io_inputs_codewords_11 : _GEN_107; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_109 = 8'hc == _GEN_32[7:0] ? io_inputs_codewords_12 : _GEN_108; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_110 = 8'hd == _GEN_32[7:0] ? io_inputs_codewords_13 : _GEN_109; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_111 = 8'he == _GEN_32[7:0] ? io_inputs_codewords_14 : _GEN_110; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_112 = 8'hf == _GEN_32[7:0] ? io_inputs_codewords_15 : _GEN_111; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_113 = 8'h10 == _GEN_32[7:0] ? io_inputs_codewords_16 : _GEN_112; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_114 = 8'h11 == _GEN_32[7:0] ? io_inputs_codewords_17 : _GEN_113; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_115 = 8'h12 == _GEN_32[7:0] ? io_inputs_codewords_18 : _GEN_114; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_116 = 8'h13 == _GEN_32[7:0] ? io_inputs_codewords_19 : _GEN_115; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_117 = 8'h14 == _GEN_32[7:0] ? io_inputs_codewords_20 : _GEN_116; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_118 = 8'h15 == _GEN_32[7:0] ? io_inputs_codewords_21 : _GEN_117; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_119 = 8'h16 == _GEN_32[7:0] ? io_inputs_codewords_22 : _GEN_118; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_120 = 8'h17 == _GEN_32[7:0] ? io_inputs_codewords_23 : _GEN_119; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_121 = 8'h18 == _GEN_32[7:0] ? io_inputs_codewords_24 : _GEN_120; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_122 = 8'h19 == _GEN_32[7:0] ? io_inputs_codewords_25 : _GEN_121; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_123 = 8'h1a == _GEN_32[7:0] ? io_inputs_codewords_26 : _GEN_122; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_124 = 8'h1b == _GEN_32[7:0] ? io_inputs_codewords_27 : _GEN_123; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_125 = 8'h1c == _GEN_32[7:0] ? io_inputs_codewords_28 : _GEN_124; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_126 = 8'h1d == _GEN_32[7:0] ? io_inputs_codewords_29 : _GEN_125; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_127 = 8'h1e == _GEN_32[7:0] ? io_inputs_codewords_30 : _GEN_126; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_128 = 8'h1f == _GEN_32[7:0] ? io_inputs_codewords_31 : _GEN_127; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_129 = 8'h20 == _GEN_32[7:0] ? io_inputs_codewords_32 : _GEN_128; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_130 = 8'h21 == _GEN_32[7:0] ? io_inputs_codewords_33 : _GEN_129; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_131 = 8'h22 == _GEN_32[7:0] ? io_inputs_codewords_34 : _GEN_130; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_132 = 8'h23 == _GEN_32[7:0] ? io_inputs_codewords_35 : _GEN_131; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_133 = 8'h24 == _GEN_32[7:0] ? io_inputs_codewords_36 : _GEN_132; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_134 = 8'h25 == _GEN_32[7:0] ? io_inputs_codewords_37 : _GEN_133; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_135 = 8'h26 == _GEN_32[7:0] ? io_inputs_codewords_38 : _GEN_134; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_136 = 8'h27 == _GEN_32[7:0] ? io_inputs_codewords_39 : _GEN_135; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_137 = 8'h28 == _GEN_32[7:0] ? io_inputs_codewords_40 : _GEN_136; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_138 = 8'h29 == _GEN_32[7:0] ? io_inputs_codewords_41 : _GEN_137; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_139 = 8'h2a == _GEN_32[7:0] ? io_inputs_codewords_42 : _GEN_138; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_140 = 8'h2b == _GEN_32[7:0] ? io_inputs_codewords_43 : _GEN_139; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_141 = 8'h2c == _GEN_32[7:0] ? io_inputs_codewords_44 : _GEN_140; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_142 = 8'h2d == _GEN_32[7:0] ? io_inputs_codewords_45 : _GEN_141; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_143 = 8'h2e == _GEN_32[7:0] ? io_inputs_codewords_46 : _GEN_142; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_144 = 8'h2f == _GEN_32[7:0] ? io_inputs_codewords_47 : _GEN_143; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_145 = 8'h30 == _GEN_32[7:0] ? io_inputs_codewords_48 : _GEN_144; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_146 = 8'h31 == _GEN_32[7:0] ? io_inputs_codewords_49 : _GEN_145; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_147 = 8'h32 == _GEN_32[7:0] ? io_inputs_codewords_50 : _GEN_146; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_148 = 8'h33 == _GEN_32[7:0] ? io_inputs_codewords_51 : _GEN_147; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_149 = 8'h34 == _GEN_32[7:0] ? io_inputs_codewords_52 : _GEN_148; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_150 = 8'h35 == _GEN_32[7:0] ? io_inputs_codewords_53 : _GEN_149; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_151 = 8'h36 == _GEN_32[7:0] ? io_inputs_codewords_54 : _GEN_150; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_152 = 8'h37 == _GEN_32[7:0] ? io_inputs_codewords_55 : _GEN_151; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_153 = 8'h38 == _GEN_32[7:0] ? io_inputs_codewords_56 : _GEN_152; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_154 = 8'h39 == _GEN_32[7:0] ? io_inputs_codewords_57 : _GEN_153; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_155 = 8'h3a == _GEN_32[7:0] ? io_inputs_codewords_58 : _GEN_154; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_156 = 8'h3b == _GEN_32[7:0] ? io_inputs_codewords_59 : _GEN_155; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_157 = 8'h3c == _GEN_32[7:0] ? io_inputs_codewords_60 : _GEN_156; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_158 = 8'h3d == _GEN_32[7:0] ? io_inputs_codewords_61 : _GEN_157; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_159 = 8'h3e == _GEN_32[7:0] ? io_inputs_codewords_62 : _GEN_158; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_160 = 8'h3f == _GEN_32[7:0] ? io_inputs_codewords_63 : _GEN_159; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_161 = 8'h40 == _GEN_32[7:0] ? io_inputs_codewords_64 : _GEN_160; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_162 = 8'h41 == _GEN_32[7:0] ? io_inputs_codewords_65 : _GEN_161; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_163 = 8'h42 == _GEN_32[7:0] ? io_inputs_codewords_66 : _GEN_162; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_164 = 8'h43 == _GEN_32[7:0] ? io_inputs_codewords_67 : _GEN_163; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_165 = 8'h44 == _GEN_32[7:0] ? io_inputs_codewords_68 : _GEN_164; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_166 = 8'h45 == _GEN_32[7:0] ? io_inputs_codewords_69 : _GEN_165; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_167 = 8'h46 == _GEN_32[7:0] ? io_inputs_codewords_70 : _GEN_166; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_168 = 8'h47 == _GEN_32[7:0] ? io_inputs_codewords_71 : _GEN_167; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_169 = 8'h48 == _GEN_32[7:0] ? io_inputs_codewords_72 : _GEN_168; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_170 = 8'h49 == _GEN_32[7:0] ? io_inputs_codewords_73 : _GEN_169; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_171 = 8'h4a == _GEN_32[7:0] ? io_inputs_codewords_74 : _GEN_170; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_172 = 8'h4b == _GEN_32[7:0] ? io_inputs_codewords_75 : _GEN_171; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_173 = 8'h4c == _GEN_32[7:0] ? io_inputs_codewords_76 : _GEN_172; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_174 = 8'h4d == _GEN_32[7:0] ? io_inputs_codewords_77 : _GEN_173; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_175 = 8'h4e == _GEN_32[7:0] ? io_inputs_codewords_78 : _GEN_174; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_176 = 8'h4f == _GEN_32[7:0] ? io_inputs_codewords_79 : _GEN_175; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_177 = 8'h50 == _GEN_32[7:0] ? io_inputs_codewords_80 : _GEN_176; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_178 = 8'h51 == _GEN_32[7:0] ? io_inputs_codewords_81 : _GEN_177; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_179 = 8'h52 == _GEN_32[7:0] ? io_inputs_codewords_82 : _GEN_178; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_180 = 8'h53 == _GEN_32[7:0] ? io_inputs_codewords_83 : _GEN_179; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_181 = 8'h54 == _GEN_32[7:0] ? io_inputs_codewords_84 : _GEN_180; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_182 = 8'h55 == _GEN_32[7:0] ? io_inputs_codewords_85 : _GEN_181; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_183 = 8'h56 == _GEN_32[7:0] ? io_inputs_codewords_86 : _GEN_182; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_184 = 8'h57 == _GEN_32[7:0] ? io_inputs_codewords_87 : _GEN_183; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_185 = 8'h58 == _GEN_32[7:0] ? io_inputs_codewords_88 : _GEN_184; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_186 = 8'h59 == _GEN_32[7:0] ? io_inputs_codewords_89 : _GEN_185; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_187 = 8'h5a == _GEN_32[7:0] ? io_inputs_codewords_90 : _GEN_186; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_188 = 8'h5b == _GEN_32[7:0] ? io_inputs_codewords_91 : _GEN_187; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_189 = 8'h5c == _GEN_32[7:0] ? io_inputs_codewords_92 : _GEN_188; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_190 = 8'h5d == _GEN_32[7:0] ? io_inputs_codewords_93 : _GEN_189; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_191 = 8'h5e == _GEN_32[7:0] ? io_inputs_codewords_94 : _GEN_190; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_192 = 8'h5f == _GEN_32[7:0] ? io_inputs_codewords_95 : _GEN_191; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_193 = 8'h60 == _GEN_32[7:0] ? io_inputs_codewords_96 : _GEN_192; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_194 = 8'h61 == _GEN_32[7:0] ? io_inputs_codewords_97 : _GEN_193; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_195 = 8'h62 == _GEN_32[7:0] ? io_inputs_codewords_98 : _GEN_194; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_196 = 8'h63 == _GEN_32[7:0] ? io_inputs_codewords_99 : _GEN_195; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_197 = 8'h64 == _GEN_32[7:0] ? io_inputs_codewords_100 : _GEN_196; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_198 = 8'h65 == _GEN_32[7:0] ? io_inputs_codewords_101 : _GEN_197; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_199 = 8'h66 == _GEN_32[7:0] ? io_inputs_codewords_102 : _GEN_198; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_200 = 8'h67 == _GEN_32[7:0] ? io_inputs_codewords_103 : _GEN_199; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_201 = 8'h68 == _GEN_32[7:0] ? io_inputs_codewords_104 : _GEN_200; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_202 = 8'h69 == _GEN_32[7:0] ? io_inputs_codewords_105 : _GEN_201; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_203 = 8'h6a == _GEN_32[7:0] ? io_inputs_codewords_106 : _GEN_202; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_204 = 8'h6b == _GEN_32[7:0] ? io_inputs_codewords_107 : _GEN_203; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_205 = 8'h6c == _GEN_32[7:0] ? io_inputs_codewords_108 : _GEN_204; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_206 = 8'h6d == _GEN_32[7:0] ? io_inputs_codewords_109 : _GEN_205; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_207 = 8'h6e == _GEN_32[7:0] ? io_inputs_codewords_110 : _GEN_206; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_208 = 8'h6f == _GEN_32[7:0] ? io_inputs_codewords_111 : _GEN_207; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_209 = 8'h70 == _GEN_32[7:0] ? io_inputs_codewords_112 : _GEN_208; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_210 = 8'h71 == _GEN_32[7:0] ? io_inputs_codewords_113 : _GEN_209; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_211 = 8'h72 == _GEN_32[7:0] ? io_inputs_codewords_114 : _GEN_210; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_212 = 8'h73 == _GEN_32[7:0] ? io_inputs_codewords_115 : _GEN_211; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_213 = 8'h74 == _GEN_32[7:0] ? io_inputs_codewords_116 : _GEN_212; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_214 = 8'h75 == _GEN_32[7:0] ? io_inputs_codewords_117 : _GEN_213; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_215 = 8'h76 == _GEN_32[7:0] ? io_inputs_codewords_118 : _GEN_214; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_216 = 8'h77 == _GEN_32[7:0] ? io_inputs_codewords_119 : _GEN_215; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_217 = 8'h78 == _GEN_32[7:0] ? io_inputs_codewords_120 : _GEN_216; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_218 = 8'h79 == _GEN_32[7:0] ? io_inputs_codewords_121 : _GEN_217; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_219 = 8'h7a == _GEN_32[7:0] ? io_inputs_codewords_122 : _GEN_218; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_220 = 8'h7b == _GEN_32[7:0] ? io_inputs_codewords_123 : _GEN_219; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_221 = 8'h7c == _GEN_32[7:0] ? io_inputs_codewords_124 : _GEN_220; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_222 = 8'h7d == _GEN_32[7:0] ? io_inputs_codewords_125 : _GEN_221; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_223 = 8'h7e == _GEN_32[7:0] ? io_inputs_codewords_126 : _GEN_222; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_224 = 8'h7f == _GEN_32[7:0] ? io_inputs_codewords_127 : _GEN_223; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_225 = 8'h80 == _GEN_32[7:0] ? io_inputs_codewords_128 : _GEN_224; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_226 = 8'h81 == _GEN_32[7:0] ? io_inputs_codewords_129 : _GEN_225; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_227 = 8'h82 == _GEN_32[7:0] ? io_inputs_codewords_130 : _GEN_226; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_228 = 8'h83 == _GEN_32[7:0] ? io_inputs_codewords_131 : _GEN_227; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_229 = 8'h84 == _GEN_32[7:0] ? io_inputs_codewords_132 : _GEN_228; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_230 = 8'h85 == _GEN_32[7:0] ? io_inputs_codewords_133 : _GEN_229; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_231 = 8'h86 == _GEN_32[7:0] ? io_inputs_codewords_134 : _GEN_230; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_232 = 8'h87 == _GEN_32[7:0] ? io_inputs_codewords_135 : _GEN_231; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_233 = 8'h88 == _GEN_32[7:0] ? io_inputs_codewords_136 : _GEN_232; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_234 = 8'h89 == _GEN_32[7:0] ? io_inputs_codewords_137 : _GEN_233; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_235 = 8'h8a == _GEN_32[7:0] ? io_inputs_codewords_138 : _GEN_234; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_236 = 8'h8b == _GEN_32[7:0] ? io_inputs_codewords_139 : _GEN_235; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_237 = 8'h8c == _GEN_32[7:0] ? io_inputs_codewords_140 : _GEN_236; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_238 = 8'h8d == _GEN_32[7:0] ? io_inputs_codewords_141 : _GEN_237; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_239 = 8'h8e == _GEN_32[7:0] ? io_inputs_codewords_142 : _GEN_238; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_240 = 8'h8f == _GEN_32[7:0] ? io_inputs_codewords_143 : _GEN_239; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_241 = 8'h90 == _GEN_32[7:0] ? io_inputs_codewords_144 : _GEN_240; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_242 = 8'h91 == _GEN_32[7:0] ? io_inputs_codewords_145 : _GEN_241; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_243 = 8'h92 == _GEN_32[7:0] ? io_inputs_codewords_146 : _GEN_242; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_244 = 8'h93 == _GEN_32[7:0] ? io_inputs_codewords_147 : _GEN_243; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_245 = 8'h94 == _GEN_32[7:0] ? io_inputs_codewords_148 : _GEN_244; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_246 = 8'h95 == _GEN_32[7:0] ? io_inputs_codewords_149 : _GEN_245; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_247 = 8'h96 == _GEN_32[7:0] ? io_inputs_codewords_150 : _GEN_246; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_248 = 8'h97 == _GEN_32[7:0] ? io_inputs_codewords_151 : _GEN_247; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_249 = 8'h98 == _GEN_32[7:0] ? io_inputs_codewords_152 : _GEN_248; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_250 = 8'h99 == _GEN_32[7:0] ? io_inputs_codewords_153 : _GEN_249; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_251 = 8'h9a == _GEN_32[7:0] ? io_inputs_codewords_154 : _GEN_250; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_252 = 8'h9b == _GEN_32[7:0] ? io_inputs_codewords_155 : _GEN_251; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_253 = 8'h9c == _GEN_32[7:0] ? io_inputs_codewords_156 : _GEN_252; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_254 = 8'h9d == _GEN_32[7:0] ? io_inputs_codewords_157 : _GEN_253; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_255 = 8'h9e == _GEN_32[7:0] ? io_inputs_codewords_158 : _GEN_254; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_256 = 8'h9f == _GEN_32[7:0] ? io_inputs_codewords_159 : _GEN_255; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_257 = 8'ha0 == _GEN_32[7:0] ? io_inputs_codewords_160 : _GEN_256; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_258 = 8'ha1 == _GEN_32[7:0] ? io_inputs_codewords_161 : _GEN_257; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_259 = 8'ha2 == _GEN_32[7:0] ? io_inputs_codewords_162 : _GEN_258; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_260 = 8'ha3 == _GEN_32[7:0] ? io_inputs_codewords_163 : _GEN_259; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_261 = 8'ha4 == _GEN_32[7:0] ? io_inputs_codewords_164 : _GEN_260; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_262 = 8'ha5 == _GEN_32[7:0] ? io_inputs_codewords_165 : _GEN_261; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_263 = 8'ha6 == _GEN_32[7:0] ? io_inputs_codewords_166 : _GEN_262; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_264 = 8'ha7 == _GEN_32[7:0] ? io_inputs_codewords_167 : _GEN_263; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_265 = 8'ha8 == _GEN_32[7:0] ? io_inputs_codewords_168 : _GEN_264; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_266 = 8'ha9 == _GEN_32[7:0] ? io_inputs_codewords_169 : _GEN_265; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_267 = 8'haa == _GEN_32[7:0] ? io_inputs_codewords_170 : _GEN_266; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_268 = 8'hab == _GEN_32[7:0] ? io_inputs_codewords_171 : _GEN_267; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_269 = 8'hac == _GEN_32[7:0] ? io_inputs_codewords_172 : _GEN_268; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_270 = 8'had == _GEN_32[7:0] ? io_inputs_codewords_173 : _GEN_269; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_271 = 8'hae == _GEN_32[7:0] ? io_inputs_codewords_174 : _GEN_270; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_272 = 8'haf == _GEN_32[7:0] ? io_inputs_codewords_175 : _GEN_271; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_273 = 8'hb0 == _GEN_32[7:0] ? io_inputs_codewords_176 : _GEN_272; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_274 = 8'hb1 == _GEN_32[7:0] ? io_inputs_codewords_177 : _GEN_273; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_275 = 8'hb2 == _GEN_32[7:0] ? io_inputs_codewords_178 : _GEN_274; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_276 = 8'hb3 == _GEN_32[7:0] ? io_inputs_codewords_179 : _GEN_275; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_277 = 8'hb4 == _GEN_32[7:0] ? io_inputs_codewords_180 : _GEN_276; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_278 = 8'hb5 == _GEN_32[7:0] ? io_inputs_codewords_181 : _GEN_277; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_279 = 8'hb6 == _GEN_32[7:0] ? io_inputs_codewords_182 : _GEN_278; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_280 = 8'hb7 == _GEN_32[7:0] ? io_inputs_codewords_183 : _GEN_279; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_281 = 8'hb8 == _GEN_32[7:0] ? io_inputs_codewords_184 : _GEN_280; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_282 = 8'hb9 == _GEN_32[7:0] ? io_inputs_codewords_185 : _GEN_281; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_283 = 8'hba == _GEN_32[7:0] ? io_inputs_codewords_186 : _GEN_282; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_284 = 8'hbb == _GEN_32[7:0] ? io_inputs_codewords_187 : _GEN_283; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_285 = 8'hbc == _GEN_32[7:0] ? io_inputs_codewords_188 : _GEN_284; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_286 = 8'hbd == _GEN_32[7:0] ? io_inputs_codewords_189 : _GEN_285; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_287 = 8'hbe == _GEN_32[7:0] ? io_inputs_codewords_190 : _GEN_286; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_288 = 8'hbf == _GEN_32[7:0] ? io_inputs_codewords_191 : _GEN_287; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_289 = 8'hc0 == _GEN_32[7:0] ? io_inputs_codewords_192 : _GEN_288; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_290 = 8'hc1 == _GEN_32[7:0] ? io_inputs_codewords_193 : _GEN_289; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_291 = 8'hc2 == _GEN_32[7:0] ? io_inputs_codewords_194 : _GEN_290; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_292 = 8'hc3 == _GEN_32[7:0] ? io_inputs_codewords_195 : _GEN_291; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_293 = 8'hc4 == _GEN_32[7:0] ? io_inputs_codewords_196 : _GEN_292; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_294 = 8'hc5 == _GEN_32[7:0] ? io_inputs_codewords_197 : _GEN_293; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_295 = 8'hc6 == _GEN_32[7:0] ? io_inputs_codewords_198 : _GEN_294; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_296 = 8'hc7 == _GEN_32[7:0] ? io_inputs_codewords_199 : _GEN_295; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_297 = 8'hc8 == _GEN_32[7:0] ? io_inputs_codewords_200 : _GEN_296; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_298 = 8'hc9 == _GEN_32[7:0] ? io_inputs_codewords_201 : _GEN_297; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_299 = 8'hca == _GEN_32[7:0] ? io_inputs_codewords_202 : _GEN_298; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_300 = 8'hcb == _GEN_32[7:0] ? io_inputs_codewords_203 : _GEN_299; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_301 = 8'hcc == _GEN_32[7:0] ? io_inputs_codewords_204 : _GEN_300; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_302 = 8'hcd == _GEN_32[7:0] ? io_inputs_codewords_205 : _GEN_301; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_303 = 8'hce == _GEN_32[7:0] ? io_inputs_codewords_206 : _GEN_302; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_304 = 8'hcf == _GEN_32[7:0] ? io_inputs_codewords_207 : _GEN_303; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_305 = 8'hd0 == _GEN_32[7:0] ? io_inputs_codewords_208 : _GEN_304; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_306 = 8'hd1 == _GEN_32[7:0] ? io_inputs_codewords_209 : _GEN_305; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_307 = 8'hd2 == _GEN_32[7:0] ? io_inputs_codewords_210 : _GEN_306; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_308 = 8'hd3 == _GEN_32[7:0] ? io_inputs_codewords_211 : _GEN_307; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_309 = 8'hd4 == _GEN_32[7:0] ? io_inputs_codewords_212 : _GEN_308; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_310 = 8'hd5 == _GEN_32[7:0] ? io_inputs_codewords_213 : _GEN_309; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_311 = 8'hd6 == _GEN_32[7:0] ? io_inputs_codewords_214 : _GEN_310; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_312 = 8'hd7 == _GEN_32[7:0] ? io_inputs_codewords_215 : _GEN_311; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_313 = 8'hd8 == _GEN_32[7:0] ? io_inputs_codewords_216 : _GEN_312; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_314 = 8'hd9 == _GEN_32[7:0] ? io_inputs_codewords_217 : _GEN_313; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_315 = 8'hda == _GEN_32[7:0] ? io_inputs_codewords_218 : _GEN_314; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_316 = 8'hdb == _GEN_32[7:0] ? io_inputs_codewords_219 : _GEN_315; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_317 = 8'hdc == _GEN_32[7:0] ? io_inputs_codewords_220 : _GEN_316; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_318 = 8'hdd == _GEN_32[7:0] ? io_inputs_codewords_221 : _GEN_317; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_319 = 8'hde == _GEN_32[7:0] ? io_inputs_codewords_222 : _GEN_318; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_320 = 8'hdf == _GEN_32[7:0] ? io_inputs_codewords_223 : _GEN_319; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_321 = 8'he0 == _GEN_32[7:0] ? io_inputs_codewords_224 : _GEN_320; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_322 = 8'he1 == _GEN_32[7:0] ? io_inputs_codewords_225 : _GEN_321; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_323 = 8'he2 == _GEN_32[7:0] ? io_inputs_codewords_226 : _GEN_322; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_324 = 8'he3 == _GEN_32[7:0] ? io_inputs_codewords_227 : _GEN_323; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_325 = 8'he4 == _GEN_32[7:0] ? io_inputs_codewords_228 : _GEN_324; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_326 = 8'he5 == _GEN_32[7:0] ? io_inputs_codewords_229 : _GEN_325; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_327 = 8'he6 == _GEN_32[7:0] ? io_inputs_codewords_230 : _GEN_326; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_328 = 8'he7 == _GEN_32[7:0] ? io_inputs_codewords_231 : _GEN_327; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_329 = 8'he8 == _GEN_32[7:0] ? io_inputs_codewords_232 : _GEN_328; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_330 = 8'he9 == _GEN_32[7:0] ? io_inputs_codewords_233 : _GEN_329; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_331 = 8'hea == _GEN_32[7:0] ? io_inputs_codewords_234 : _GEN_330; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_332 = 8'heb == _GEN_32[7:0] ? io_inputs_codewords_235 : _GEN_331; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_333 = 8'hec == _GEN_32[7:0] ? io_inputs_codewords_236 : _GEN_332; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_334 = 8'hed == _GEN_32[7:0] ? io_inputs_codewords_237 : _GEN_333; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_335 = 8'hee == _GEN_32[7:0] ? io_inputs_codewords_238 : _GEN_334; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_336 = 8'hef == _GEN_32[7:0] ? io_inputs_codewords_239 : _GEN_335; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_337 = 8'hf0 == _GEN_32[7:0] ? io_inputs_codewords_240 : _GEN_336; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_338 = 8'hf1 == _GEN_32[7:0] ? io_inputs_codewords_241 : _GEN_337; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_339 = 8'hf2 == _GEN_32[7:0] ? io_inputs_codewords_242 : _GEN_338; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_340 = 8'hf3 == _GEN_32[7:0] ? io_inputs_codewords_243 : _GEN_339; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_341 = 8'hf4 == _GEN_32[7:0] ? io_inputs_codewords_244 : _GEN_340; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_342 = 8'hf5 == _GEN_32[7:0] ? io_inputs_codewords_245 : _GEN_341; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_343 = 8'hf6 == _GEN_32[7:0] ? io_inputs_codewords_246 : _GEN_342; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_344 = 8'hf7 == _GEN_32[7:0] ? io_inputs_codewords_247 : _GEN_343; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_345 = 8'hf8 == _GEN_32[7:0] ? io_inputs_codewords_248 : _GEN_344; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_346 = 8'hf9 == _GEN_32[7:0] ? io_inputs_codewords_249 : _GEN_345; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_347 = 8'hfa == _GEN_32[7:0] ? io_inputs_codewords_250 : _GEN_346; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_348 = 8'hfb == _GEN_32[7:0] ? io_inputs_codewords_251 : _GEN_347; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_349 = 8'hfc == _GEN_32[7:0] ? io_inputs_codewords_252 : _GEN_348; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_350 = 8'hfd == _GEN_32[7:0] ? io_inputs_codewords_253 : _GEN_349; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_351 = 8'hfe == _GEN_32[7:0] ? io_inputs_codewords_254 : _GEN_350; // @[compressorOutput.scala 104:74]
  wire [23:0] _GEN_352 = 8'hff == _GEN_32[7:0] ? io_inputs_codewords_255 : _GEN_351; // @[compressorOutput.scala 104:74]
  wire [4:0] _GEN_386 = 8'h1 == _GEN_32[7:0] ? io_inputs_lengths_1 : io_inputs_lengths_0; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_387 = 8'h2 == _GEN_32[7:0] ? io_inputs_lengths_2 : _GEN_386; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_388 = 8'h3 == _GEN_32[7:0] ? io_inputs_lengths_3 : _GEN_387; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_389 = 8'h4 == _GEN_32[7:0] ? io_inputs_lengths_4 : _GEN_388; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_390 = 8'h5 == _GEN_32[7:0] ? io_inputs_lengths_5 : _GEN_389; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_391 = 8'h6 == _GEN_32[7:0] ? io_inputs_lengths_6 : _GEN_390; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_392 = 8'h7 == _GEN_32[7:0] ? io_inputs_lengths_7 : _GEN_391; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_393 = 8'h8 == _GEN_32[7:0] ? io_inputs_lengths_8 : _GEN_392; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_394 = 8'h9 == _GEN_32[7:0] ? io_inputs_lengths_9 : _GEN_393; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_395 = 8'ha == _GEN_32[7:0] ? io_inputs_lengths_10 : _GEN_394; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_396 = 8'hb == _GEN_32[7:0] ? io_inputs_lengths_11 : _GEN_395; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_397 = 8'hc == _GEN_32[7:0] ? io_inputs_lengths_12 : _GEN_396; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_398 = 8'hd == _GEN_32[7:0] ? io_inputs_lengths_13 : _GEN_397; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_399 = 8'he == _GEN_32[7:0] ? io_inputs_lengths_14 : _GEN_398; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_400 = 8'hf == _GEN_32[7:0] ? io_inputs_lengths_15 : _GEN_399; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_401 = 8'h10 == _GEN_32[7:0] ? io_inputs_lengths_16 : _GEN_400; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_402 = 8'h11 == _GEN_32[7:0] ? io_inputs_lengths_17 : _GEN_401; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_403 = 8'h12 == _GEN_32[7:0] ? io_inputs_lengths_18 : _GEN_402; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_404 = 8'h13 == _GEN_32[7:0] ? io_inputs_lengths_19 : _GEN_403; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_405 = 8'h14 == _GEN_32[7:0] ? io_inputs_lengths_20 : _GEN_404; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_406 = 8'h15 == _GEN_32[7:0] ? io_inputs_lengths_21 : _GEN_405; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_407 = 8'h16 == _GEN_32[7:0] ? io_inputs_lengths_22 : _GEN_406; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_408 = 8'h17 == _GEN_32[7:0] ? io_inputs_lengths_23 : _GEN_407; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_409 = 8'h18 == _GEN_32[7:0] ? io_inputs_lengths_24 : _GEN_408; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_410 = 8'h19 == _GEN_32[7:0] ? io_inputs_lengths_25 : _GEN_409; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_411 = 8'h1a == _GEN_32[7:0] ? io_inputs_lengths_26 : _GEN_410; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_412 = 8'h1b == _GEN_32[7:0] ? io_inputs_lengths_27 : _GEN_411; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_413 = 8'h1c == _GEN_32[7:0] ? io_inputs_lengths_28 : _GEN_412; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_414 = 8'h1d == _GEN_32[7:0] ? io_inputs_lengths_29 : _GEN_413; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_415 = 8'h1e == _GEN_32[7:0] ? io_inputs_lengths_30 : _GEN_414; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_416 = 8'h1f == _GEN_32[7:0] ? io_inputs_lengths_31 : _GEN_415; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_417 = 8'h20 == _GEN_32[7:0] ? io_inputs_lengths_32 : _GEN_416; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_418 = 8'h21 == _GEN_32[7:0] ? io_inputs_lengths_33 : _GEN_417; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_419 = 8'h22 == _GEN_32[7:0] ? io_inputs_lengths_34 : _GEN_418; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_420 = 8'h23 == _GEN_32[7:0] ? io_inputs_lengths_35 : _GEN_419; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_421 = 8'h24 == _GEN_32[7:0] ? io_inputs_lengths_36 : _GEN_420; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_422 = 8'h25 == _GEN_32[7:0] ? io_inputs_lengths_37 : _GEN_421; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_423 = 8'h26 == _GEN_32[7:0] ? io_inputs_lengths_38 : _GEN_422; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_424 = 8'h27 == _GEN_32[7:0] ? io_inputs_lengths_39 : _GEN_423; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_425 = 8'h28 == _GEN_32[7:0] ? io_inputs_lengths_40 : _GEN_424; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_426 = 8'h29 == _GEN_32[7:0] ? io_inputs_lengths_41 : _GEN_425; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_427 = 8'h2a == _GEN_32[7:0] ? io_inputs_lengths_42 : _GEN_426; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_428 = 8'h2b == _GEN_32[7:0] ? io_inputs_lengths_43 : _GEN_427; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_429 = 8'h2c == _GEN_32[7:0] ? io_inputs_lengths_44 : _GEN_428; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_430 = 8'h2d == _GEN_32[7:0] ? io_inputs_lengths_45 : _GEN_429; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_431 = 8'h2e == _GEN_32[7:0] ? io_inputs_lengths_46 : _GEN_430; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_432 = 8'h2f == _GEN_32[7:0] ? io_inputs_lengths_47 : _GEN_431; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_433 = 8'h30 == _GEN_32[7:0] ? io_inputs_lengths_48 : _GEN_432; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_434 = 8'h31 == _GEN_32[7:0] ? io_inputs_lengths_49 : _GEN_433; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_435 = 8'h32 == _GEN_32[7:0] ? io_inputs_lengths_50 : _GEN_434; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_436 = 8'h33 == _GEN_32[7:0] ? io_inputs_lengths_51 : _GEN_435; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_437 = 8'h34 == _GEN_32[7:0] ? io_inputs_lengths_52 : _GEN_436; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_438 = 8'h35 == _GEN_32[7:0] ? io_inputs_lengths_53 : _GEN_437; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_439 = 8'h36 == _GEN_32[7:0] ? io_inputs_lengths_54 : _GEN_438; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_440 = 8'h37 == _GEN_32[7:0] ? io_inputs_lengths_55 : _GEN_439; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_441 = 8'h38 == _GEN_32[7:0] ? io_inputs_lengths_56 : _GEN_440; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_442 = 8'h39 == _GEN_32[7:0] ? io_inputs_lengths_57 : _GEN_441; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_443 = 8'h3a == _GEN_32[7:0] ? io_inputs_lengths_58 : _GEN_442; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_444 = 8'h3b == _GEN_32[7:0] ? io_inputs_lengths_59 : _GEN_443; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_445 = 8'h3c == _GEN_32[7:0] ? io_inputs_lengths_60 : _GEN_444; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_446 = 8'h3d == _GEN_32[7:0] ? io_inputs_lengths_61 : _GEN_445; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_447 = 8'h3e == _GEN_32[7:0] ? io_inputs_lengths_62 : _GEN_446; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_448 = 8'h3f == _GEN_32[7:0] ? io_inputs_lengths_63 : _GEN_447; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_449 = 8'h40 == _GEN_32[7:0] ? io_inputs_lengths_64 : _GEN_448; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_450 = 8'h41 == _GEN_32[7:0] ? io_inputs_lengths_65 : _GEN_449; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_451 = 8'h42 == _GEN_32[7:0] ? io_inputs_lengths_66 : _GEN_450; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_452 = 8'h43 == _GEN_32[7:0] ? io_inputs_lengths_67 : _GEN_451; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_453 = 8'h44 == _GEN_32[7:0] ? io_inputs_lengths_68 : _GEN_452; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_454 = 8'h45 == _GEN_32[7:0] ? io_inputs_lengths_69 : _GEN_453; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_455 = 8'h46 == _GEN_32[7:0] ? io_inputs_lengths_70 : _GEN_454; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_456 = 8'h47 == _GEN_32[7:0] ? io_inputs_lengths_71 : _GEN_455; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_457 = 8'h48 == _GEN_32[7:0] ? io_inputs_lengths_72 : _GEN_456; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_458 = 8'h49 == _GEN_32[7:0] ? io_inputs_lengths_73 : _GEN_457; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_459 = 8'h4a == _GEN_32[7:0] ? io_inputs_lengths_74 : _GEN_458; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_460 = 8'h4b == _GEN_32[7:0] ? io_inputs_lengths_75 : _GEN_459; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_461 = 8'h4c == _GEN_32[7:0] ? io_inputs_lengths_76 : _GEN_460; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_462 = 8'h4d == _GEN_32[7:0] ? io_inputs_lengths_77 : _GEN_461; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_463 = 8'h4e == _GEN_32[7:0] ? io_inputs_lengths_78 : _GEN_462; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_464 = 8'h4f == _GEN_32[7:0] ? io_inputs_lengths_79 : _GEN_463; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_465 = 8'h50 == _GEN_32[7:0] ? io_inputs_lengths_80 : _GEN_464; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_466 = 8'h51 == _GEN_32[7:0] ? io_inputs_lengths_81 : _GEN_465; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_467 = 8'h52 == _GEN_32[7:0] ? io_inputs_lengths_82 : _GEN_466; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_468 = 8'h53 == _GEN_32[7:0] ? io_inputs_lengths_83 : _GEN_467; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_469 = 8'h54 == _GEN_32[7:0] ? io_inputs_lengths_84 : _GEN_468; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_470 = 8'h55 == _GEN_32[7:0] ? io_inputs_lengths_85 : _GEN_469; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_471 = 8'h56 == _GEN_32[7:0] ? io_inputs_lengths_86 : _GEN_470; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_472 = 8'h57 == _GEN_32[7:0] ? io_inputs_lengths_87 : _GEN_471; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_473 = 8'h58 == _GEN_32[7:0] ? io_inputs_lengths_88 : _GEN_472; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_474 = 8'h59 == _GEN_32[7:0] ? io_inputs_lengths_89 : _GEN_473; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_475 = 8'h5a == _GEN_32[7:0] ? io_inputs_lengths_90 : _GEN_474; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_476 = 8'h5b == _GEN_32[7:0] ? io_inputs_lengths_91 : _GEN_475; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_477 = 8'h5c == _GEN_32[7:0] ? io_inputs_lengths_92 : _GEN_476; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_478 = 8'h5d == _GEN_32[7:0] ? io_inputs_lengths_93 : _GEN_477; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_479 = 8'h5e == _GEN_32[7:0] ? io_inputs_lengths_94 : _GEN_478; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_480 = 8'h5f == _GEN_32[7:0] ? io_inputs_lengths_95 : _GEN_479; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_481 = 8'h60 == _GEN_32[7:0] ? io_inputs_lengths_96 : _GEN_480; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_482 = 8'h61 == _GEN_32[7:0] ? io_inputs_lengths_97 : _GEN_481; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_483 = 8'h62 == _GEN_32[7:0] ? io_inputs_lengths_98 : _GEN_482; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_484 = 8'h63 == _GEN_32[7:0] ? io_inputs_lengths_99 : _GEN_483; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_485 = 8'h64 == _GEN_32[7:0] ? io_inputs_lengths_100 : _GEN_484; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_486 = 8'h65 == _GEN_32[7:0] ? io_inputs_lengths_101 : _GEN_485; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_487 = 8'h66 == _GEN_32[7:0] ? io_inputs_lengths_102 : _GEN_486; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_488 = 8'h67 == _GEN_32[7:0] ? io_inputs_lengths_103 : _GEN_487; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_489 = 8'h68 == _GEN_32[7:0] ? io_inputs_lengths_104 : _GEN_488; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_490 = 8'h69 == _GEN_32[7:0] ? io_inputs_lengths_105 : _GEN_489; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_491 = 8'h6a == _GEN_32[7:0] ? io_inputs_lengths_106 : _GEN_490; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_492 = 8'h6b == _GEN_32[7:0] ? io_inputs_lengths_107 : _GEN_491; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_493 = 8'h6c == _GEN_32[7:0] ? io_inputs_lengths_108 : _GEN_492; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_494 = 8'h6d == _GEN_32[7:0] ? io_inputs_lengths_109 : _GEN_493; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_495 = 8'h6e == _GEN_32[7:0] ? io_inputs_lengths_110 : _GEN_494; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_496 = 8'h6f == _GEN_32[7:0] ? io_inputs_lengths_111 : _GEN_495; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_497 = 8'h70 == _GEN_32[7:0] ? io_inputs_lengths_112 : _GEN_496; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_498 = 8'h71 == _GEN_32[7:0] ? io_inputs_lengths_113 : _GEN_497; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_499 = 8'h72 == _GEN_32[7:0] ? io_inputs_lengths_114 : _GEN_498; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_500 = 8'h73 == _GEN_32[7:0] ? io_inputs_lengths_115 : _GEN_499; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_501 = 8'h74 == _GEN_32[7:0] ? io_inputs_lengths_116 : _GEN_500; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_502 = 8'h75 == _GEN_32[7:0] ? io_inputs_lengths_117 : _GEN_501; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_503 = 8'h76 == _GEN_32[7:0] ? io_inputs_lengths_118 : _GEN_502; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_504 = 8'h77 == _GEN_32[7:0] ? io_inputs_lengths_119 : _GEN_503; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_505 = 8'h78 == _GEN_32[7:0] ? io_inputs_lengths_120 : _GEN_504; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_506 = 8'h79 == _GEN_32[7:0] ? io_inputs_lengths_121 : _GEN_505; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_507 = 8'h7a == _GEN_32[7:0] ? io_inputs_lengths_122 : _GEN_506; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_508 = 8'h7b == _GEN_32[7:0] ? io_inputs_lengths_123 : _GEN_507; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_509 = 8'h7c == _GEN_32[7:0] ? io_inputs_lengths_124 : _GEN_508; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_510 = 8'h7d == _GEN_32[7:0] ? io_inputs_lengths_125 : _GEN_509; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_511 = 8'h7e == _GEN_32[7:0] ? io_inputs_lengths_126 : _GEN_510; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_512 = 8'h7f == _GEN_32[7:0] ? io_inputs_lengths_127 : _GEN_511; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_513 = 8'h80 == _GEN_32[7:0] ? io_inputs_lengths_128 : _GEN_512; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_514 = 8'h81 == _GEN_32[7:0] ? io_inputs_lengths_129 : _GEN_513; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_515 = 8'h82 == _GEN_32[7:0] ? io_inputs_lengths_130 : _GEN_514; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_516 = 8'h83 == _GEN_32[7:0] ? io_inputs_lengths_131 : _GEN_515; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_517 = 8'h84 == _GEN_32[7:0] ? io_inputs_lengths_132 : _GEN_516; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_518 = 8'h85 == _GEN_32[7:0] ? io_inputs_lengths_133 : _GEN_517; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_519 = 8'h86 == _GEN_32[7:0] ? io_inputs_lengths_134 : _GEN_518; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_520 = 8'h87 == _GEN_32[7:0] ? io_inputs_lengths_135 : _GEN_519; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_521 = 8'h88 == _GEN_32[7:0] ? io_inputs_lengths_136 : _GEN_520; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_522 = 8'h89 == _GEN_32[7:0] ? io_inputs_lengths_137 : _GEN_521; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_523 = 8'h8a == _GEN_32[7:0] ? io_inputs_lengths_138 : _GEN_522; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_524 = 8'h8b == _GEN_32[7:0] ? io_inputs_lengths_139 : _GEN_523; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_525 = 8'h8c == _GEN_32[7:0] ? io_inputs_lengths_140 : _GEN_524; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_526 = 8'h8d == _GEN_32[7:0] ? io_inputs_lengths_141 : _GEN_525; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_527 = 8'h8e == _GEN_32[7:0] ? io_inputs_lengths_142 : _GEN_526; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_528 = 8'h8f == _GEN_32[7:0] ? io_inputs_lengths_143 : _GEN_527; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_529 = 8'h90 == _GEN_32[7:0] ? io_inputs_lengths_144 : _GEN_528; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_530 = 8'h91 == _GEN_32[7:0] ? io_inputs_lengths_145 : _GEN_529; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_531 = 8'h92 == _GEN_32[7:0] ? io_inputs_lengths_146 : _GEN_530; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_532 = 8'h93 == _GEN_32[7:0] ? io_inputs_lengths_147 : _GEN_531; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_533 = 8'h94 == _GEN_32[7:0] ? io_inputs_lengths_148 : _GEN_532; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_534 = 8'h95 == _GEN_32[7:0] ? io_inputs_lengths_149 : _GEN_533; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_535 = 8'h96 == _GEN_32[7:0] ? io_inputs_lengths_150 : _GEN_534; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_536 = 8'h97 == _GEN_32[7:0] ? io_inputs_lengths_151 : _GEN_535; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_537 = 8'h98 == _GEN_32[7:0] ? io_inputs_lengths_152 : _GEN_536; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_538 = 8'h99 == _GEN_32[7:0] ? io_inputs_lengths_153 : _GEN_537; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_539 = 8'h9a == _GEN_32[7:0] ? io_inputs_lengths_154 : _GEN_538; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_540 = 8'h9b == _GEN_32[7:0] ? io_inputs_lengths_155 : _GEN_539; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_541 = 8'h9c == _GEN_32[7:0] ? io_inputs_lengths_156 : _GEN_540; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_542 = 8'h9d == _GEN_32[7:0] ? io_inputs_lengths_157 : _GEN_541; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_543 = 8'h9e == _GEN_32[7:0] ? io_inputs_lengths_158 : _GEN_542; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_544 = 8'h9f == _GEN_32[7:0] ? io_inputs_lengths_159 : _GEN_543; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_545 = 8'ha0 == _GEN_32[7:0] ? io_inputs_lengths_160 : _GEN_544; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_546 = 8'ha1 == _GEN_32[7:0] ? io_inputs_lengths_161 : _GEN_545; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_547 = 8'ha2 == _GEN_32[7:0] ? io_inputs_lengths_162 : _GEN_546; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_548 = 8'ha3 == _GEN_32[7:0] ? io_inputs_lengths_163 : _GEN_547; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_549 = 8'ha4 == _GEN_32[7:0] ? io_inputs_lengths_164 : _GEN_548; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_550 = 8'ha5 == _GEN_32[7:0] ? io_inputs_lengths_165 : _GEN_549; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_551 = 8'ha6 == _GEN_32[7:0] ? io_inputs_lengths_166 : _GEN_550; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_552 = 8'ha7 == _GEN_32[7:0] ? io_inputs_lengths_167 : _GEN_551; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_553 = 8'ha8 == _GEN_32[7:0] ? io_inputs_lengths_168 : _GEN_552; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_554 = 8'ha9 == _GEN_32[7:0] ? io_inputs_lengths_169 : _GEN_553; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_555 = 8'haa == _GEN_32[7:0] ? io_inputs_lengths_170 : _GEN_554; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_556 = 8'hab == _GEN_32[7:0] ? io_inputs_lengths_171 : _GEN_555; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_557 = 8'hac == _GEN_32[7:0] ? io_inputs_lengths_172 : _GEN_556; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_558 = 8'had == _GEN_32[7:0] ? io_inputs_lengths_173 : _GEN_557; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_559 = 8'hae == _GEN_32[7:0] ? io_inputs_lengths_174 : _GEN_558; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_560 = 8'haf == _GEN_32[7:0] ? io_inputs_lengths_175 : _GEN_559; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_561 = 8'hb0 == _GEN_32[7:0] ? io_inputs_lengths_176 : _GEN_560; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_562 = 8'hb1 == _GEN_32[7:0] ? io_inputs_lengths_177 : _GEN_561; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_563 = 8'hb2 == _GEN_32[7:0] ? io_inputs_lengths_178 : _GEN_562; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_564 = 8'hb3 == _GEN_32[7:0] ? io_inputs_lengths_179 : _GEN_563; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_565 = 8'hb4 == _GEN_32[7:0] ? io_inputs_lengths_180 : _GEN_564; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_566 = 8'hb5 == _GEN_32[7:0] ? io_inputs_lengths_181 : _GEN_565; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_567 = 8'hb6 == _GEN_32[7:0] ? io_inputs_lengths_182 : _GEN_566; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_568 = 8'hb7 == _GEN_32[7:0] ? io_inputs_lengths_183 : _GEN_567; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_569 = 8'hb8 == _GEN_32[7:0] ? io_inputs_lengths_184 : _GEN_568; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_570 = 8'hb9 == _GEN_32[7:0] ? io_inputs_lengths_185 : _GEN_569; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_571 = 8'hba == _GEN_32[7:0] ? io_inputs_lengths_186 : _GEN_570; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_572 = 8'hbb == _GEN_32[7:0] ? io_inputs_lengths_187 : _GEN_571; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_573 = 8'hbc == _GEN_32[7:0] ? io_inputs_lengths_188 : _GEN_572; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_574 = 8'hbd == _GEN_32[7:0] ? io_inputs_lengths_189 : _GEN_573; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_575 = 8'hbe == _GEN_32[7:0] ? io_inputs_lengths_190 : _GEN_574; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_576 = 8'hbf == _GEN_32[7:0] ? io_inputs_lengths_191 : _GEN_575; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_577 = 8'hc0 == _GEN_32[7:0] ? io_inputs_lengths_192 : _GEN_576; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_578 = 8'hc1 == _GEN_32[7:0] ? io_inputs_lengths_193 : _GEN_577; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_579 = 8'hc2 == _GEN_32[7:0] ? io_inputs_lengths_194 : _GEN_578; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_580 = 8'hc3 == _GEN_32[7:0] ? io_inputs_lengths_195 : _GEN_579; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_581 = 8'hc4 == _GEN_32[7:0] ? io_inputs_lengths_196 : _GEN_580; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_582 = 8'hc5 == _GEN_32[7:0] ? io_inputs_lengths_197 : _GEN_581; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_583 = 8'hc6 == _GEN_32[7:0] ? io_inputs_lengths_198 : _GEN_582; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_584 = 8'hc7 == _GEN_32[7:0] ? io_inputs_lengths_199 : _GEN_583; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_585 = 8'hc8 == _GEN_32[7:0] ? io_inputs_lengths_200 : _GEN_584; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_586 = 8'hc9 == _GEN_32[7:0] ? io_inputs_lengths_201 : _GEN_585; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_587 = 8'hca == _GEN_32[7:0] ? io_inputs_lengths_202 : _GEN_586; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_588 = 8'hcb == _GEN_32[7:0] ? io_inputs_lengths_203 : _GEN_587; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_589 = 8'hcc == _GEN_32[7:0] ? io_inputs_lengths_204 : _GEN_588; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_590 = 8'hcd == _GEN_32[7:0] ? io_inputs_lengths_205 : _GEN_589; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_591 = 8'hce == _GEN_32[7:0] ? io_inputs_lengths_206 : _GEN_590; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_592 = 8'hcf == _GEN_32[7:0] ? io_inputs_lengths_207 : _GEN_591; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_593 = 8'hd0 == _GEN_32[7:0] ? io_inputs_lengths_208 : _GEN_592; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_594 = 8'hd1 == _GEN_32[7:0] ? io_inputs_lengths_209 : _GEN_593; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_595 = 8'hd2 == _GEN_32[7:0] ? io_inputs_lengths_210 : _GEN_594; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_596 = 8'hd3 == _GEN_32[7:0] ? io_inputs_lengths_211 : _GEN_595; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_597 = 8'hd4 == _GEN_32[7:0] ? io_inputs_lengths_212 : _GEN_596; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_598 = 8'hd5 == _GEN_32[7:0] ? io_inputs_lengths_213 : _GEN_597; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_599 = 8'hd6 == _GEN_32[7:0] ? io_inputs_lengths_214 : _GEN_598; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_600 = 8'hd7 == _GEN_32[7:0] ? io_inputs_lengths_215 : _GEN_599; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_601 = 8'hd8 == _GEN_32[7:0] ? io_inputs_lengths_216 : _GEN_600; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_602 = 8'hd9 == _GEN_32[7:0] ? io_inputs_lengths_217 : _GEN_601; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_603 = 8'hda == _GEN_32[7:0] ? io_inputs_lengths_218 : _GEN_602; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_604 = 8'hdb == _GEN_32[7:0] ? io_inputs_lengths_219 : _GEN_603; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_605 = 8'hdc == _GEN_32[7:0] ? io_inputs_lengths_220 : _GEN_604; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_606 = 8'hdd == _GEN_32[7:0] ? io_inputs_lengths_221 : _GEN_605; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_607 = 8'hde == _GEN_32[7:0] ? io_inputs_lengths_222 : _GEN_606; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_608 = 8'hdf == _GEN_32[7:0] ? io_inputs_lengths_223 : _GEN_607; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_609 = 8'he0 == _GEN_32[7:0] ? io_inputs_lengths_224 : _GEN_608; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_610 = 8'he1 == _GEN_32[7:0] ? io_inputs_lengths_225 : _GEN_609; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_611 = 8'he2 == _GEN_32[7:0] ? io_inputs_lengths_226 : _GEN_610; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_612 = 8'he3 == _GEN_32[7:0] ? io_inputs_lengths_227 : _GEN_611; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_613 = 8'he4 == _GEN_32[7:0] ? io_inputs_lengths_228 : _GEN_612; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_614 = 8'he5 == _GEN_32[7:0] ? io_inputs_lengths_229 : _GEN_613; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_615 = 8'he6 == _GEN_32[7:0] ? io_inputs_lengths_230 : _GEN_614; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_616 = 8'he7 == _GEN_32[7:0] ? io_inputs_lengths_231 : _GEN_615; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_617 = 8'he8 == _GEN_32[7:0] ? io_inputs_lengths_232 : _GEN_616; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_618 = 8'he9 == _GEN_32[7:0] ? io_inputs_lengths_233 : _GEN_617; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_619 = 8'hea == _GEN_32[7:0] ? io_inputs_lengths_234 : _GEN_618; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_620 = 8'heb == _GEN_32[7:0] ? io_inputs_lengths_235 : _GEN_619; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_621 = 8'hec == _GEN_32[7:0] ? io_inputs_lengths_236 : _GEN_620; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_622 = 8'hed == _GEN_32[7:0] ? io_inputs_lengths_237 : _GEN_621; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_623 = 8'hee == _GEN_32[7:0] ? io_inputs_lengths_238 : _GEN_622; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_624 = 8'hef == _GEN_32[7:0] ? io_inputs_lengths_239 : _GEN_623; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_625 = 8'hf0 == _GEN_32[7:0] ? io_inputs_lengths_240 : _GEN_624; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_626 = 8'hf1 == _GEN_32[7:0] ? io_inputs_lengths_241 : _GEN_625; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_627 = 8'hf2 == _GEN_32[7:0] ? io_inputs_lengths_242 : _GEN_626; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_628 = 8'hf3 == _GEN_32[7:0] ? io_inputs_lengths_243 : _GEN_627; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_629 = 8'hf4 == _GEN_32[7:0] ? io_inputs_lengths_244 : _GEN_628; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_630 = 8'hf5 == _GEN_32[7:0] ? io_inputs_lengths_245 : _GEN_629; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_631 = 8'hf6 == _GEN_32[7:0] ? io_inputs_lengths_246 : _GEN_630; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_632 = 8'hf7 == _GEN_32[7:0] ? io_inputs_lengths_247 : _GEN_631; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_633 = 8'hf8 == _GEN_32[7:0] ? io_inputs_lengths_248 : _GEN_632; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_634 = 8'hf9 == _GEN_32[7:0] ? io_inputs_lengths_249 : _GEN_633; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_635 = 8'hfa == _GEN_32[7:0] ? io_inputs_lengths_250 : _GEN_634; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_636 = 8'hfb == _GEN_32[7:0] ? io_inputs_lengths_251 : _GEN_635; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_637 = 8'hfc == _GEN_32[7:0] ? io_inputs_lengths_252 : _GEN_636; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_638 = 8'hfd == _GEN_32[7:0] ? io_inputs_lengths_253 : _GEN_637; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_639 = 8'hfe == _GEN_32[7:0] ? io_inputs_lengths_254 : _GEN_638; // @[compressorOutput.scala 108:72]
  wire [4:0] _GEN_640 = 8'hff == _GEN_32[7:0] ? io_inputs_lengths_255 : _GEN_639; // @[compressorOutput.scala 108:72]
  wire [27:0] _T_18 = {_GEN_32,_GEN_352[14:0],_GEN_640[3:0]}; // @[Cat.scala 29:58]
  wire [27:0] _GEN_673 = _GEN_32[8] ? _T_9 : _T_18; // @[compressorOutput.scala 90:11]
  wire [27:0] _GEN_674 = _T_2 ? _GEN_673 : 28'h0; // @[compressorOutput.scala 87:45]
  wire [12:0] _T_20 = iterations_0 + 13'h1; // @[compressorOutput.scala 121:40]
  wire  _T_23 = _T_20 >= 13'h20; // @[compressorOutput.scala 122:34]
  wire  _T_24 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_25 = iterations_0 < 13'h1000; // @[compressorOutput.scala 135:60]
  wire [13:0] _T_26 = {{1'd0}, iterations_0}; // @[compressorOutput.scala 136:58]
  wire [4:0] _GEN_680 = 8'h1 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_1 : io_inputs_lengths_0; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_681 = 8'h2 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_2 : _GEN_680; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_682 = 8'h3 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_3 : _GEN_681; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_683 = 8'h4 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_4 : _GEN_682; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_684 = 8'h5 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_5 : _GEN_683; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_685 = 8'h6 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_6 : _GEN_684; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_686 = 8'h7 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_7 : _GEN_685; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_687 = 8'h8 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_8 : _GEN_686; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_688 = 8'h9 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_9 : _GEN_687; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_689 = 8'ha == input_0_io_dataOut_bits_0 ? io_inputs_lengths_10 : _GEN_688; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_690 = 8'hb == input_0_io_dataOut_bits_0 ? io_inputs_lengths_11 : _GEN_689; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_691 = 8'hc == input_0_io_dataOut_bits_0 ? io_inputs_lengths_12 : _GEN_690; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_692 = 8'hd == input_0_io_dataOut_bits_0 ? io_inputs_lengths_13 : _GEN_691; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_693 = 8'he == input_0_io_dataOut_bits_0 ? io_inputs_lengths_14 : _GEN_692; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_694 = 8'hf == input_0_io_dataOut_bits_0 ? io_inputs_lengths_15 : _GEN_693; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_695 = 8'h10 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_16 : _GEN_694; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_696 = 8'h11 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_17 : _GEN_695; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_697 = 8'h12 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_18 : _GEN_696; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_698 = 8'h13 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_19 : _GEN_697; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_699 = 8'h14 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_20 : _GEN_698; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_700 = 8'h15 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_21 : _GEN_699; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_701 = 8'h16 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_22 : _GEN_700; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_702 = 8'h17 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_23 : _GEN_701; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_703 = 8'h18 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_24 : _GEN_702; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_704 = 8'h19 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_25 : _GEN_703; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_705 = 8'h1a == input_0_io_dataOut_bits_0 ? io_inputs_lengths_26 : _GEN_704; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_706 = 8'h1b == input_0_io_dataOut_bits_0 ? io_inputs_lengths_27 : _GEN_705; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_707 = 8'h1c == input_0_io_dataOut_bits_0 ? io_inputs_lengths_28 : _GEN_706; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_708 = 8'h1d == input_0_io_dataOut_bits_0 ? io_inputs_lengths_29 : _GEN_707; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_709 = 8'h1e == input_0_io_dataOut_bits_0 ? io_inputs_lengths_30 : _GEN_708; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_710 = 8'h1f == input_0_io_dataOut_bits_0 ? io_inputs_lengths_31 : _GEN_709; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_711 = 8'h20 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_32 : _GEN_710; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_712 = 8'h21 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_33 : _GEN_711; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_713 = 8'h22 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_34 : _GEN_712; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_714 = 8'h23 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_35 : _GEN_713; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_715 = 8'h24 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_36 : _GEN_714; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_716 = 8'h25 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_37 : _GEN_715; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_717 = 8'h26 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_38 : _GEN_716; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_718 = 8'h27 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_39 : _GEN_717; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_719 = 8'h28 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_40 : _GEN_718; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_720 = 8'h29 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_41 : _GEN_719; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_721 = 8'h2a == input_0_io_dataOut_bits_0 ? io_inputs_lengths_42 : _GEN_720; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_722 = 8'h2b == input_0_io_dataOut_bits_0 ? io_inputs_lengths_43 : _GEN_721; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_723 = 8'h2c == input_0_io_dataOut_bits_0 ? io_inputs_lengths_44 : _GEN_722; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_724 = 8'h2d == input_0_io_dataOut_bits_0 ? io_inputs_lengths_45 : _GEN_723; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_725 = 8'h2e == input_0_io_dataOut_bits_0 ? io_inputs_lengths_46 : _GEN_724; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_726 = 8'h2f == input_0_io_dataOut_bits_0 ? io_inputs_lengths_47 : _GEN_725; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_727 = 8'h30 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_48 : _GEN_726; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_728 = 8'h31 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_49 : _GEN_727; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_729 = 8'h32 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_50 : _GEN_728; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_730 = 8'h33 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_51 : _GEN_729; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_731 = 8'h34 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_52 : _GEN_730; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_732 = 8'h35 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_53 : _GEN_731; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_733 = 8'h36 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_54 : _GEN_732; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_734 = 8'h37 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_55 : _GEN_733; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_735 = 8'h38 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_56 : _GEN_734; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_736 = 8'h39 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_57 : _GEN_735; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_737 = 8'h3a == input_0_io_dataOut_bits_0 ? io_inputs_lengths_58 : _GEN_736; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_738 = 8'h3b == input_0_io_dataOut_bits_0 ? io_inputs_lengths_59 : _GEN_737; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_739 = 8'h3c == input_0_io_dataOut_bits_0 ? io_inputs_lengths_60 : _GEN_738; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_740 = 8'h3d == input_0_io_dataOut_bits_0 ? io_inputs_lengths_61 : _GEN_739; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_741 = 8'h3e == input_0_io_dataOut_bits_0 ? io_inputs_lengths_62 : _GEN_740; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_742 = 8'h3f == input_0_io_dataOut_bits_0 ? io_inputs_lengths_63 : _GEN_741; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_743 = 8'h40 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_64 : _GEN_742; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_744 = 8'h41 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_65 : _GEN_743; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_745 = 8'h42 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_66 : _GEN_744; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_746 = 8'h43 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_67 : _GEN_745; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_747 = 8'h44 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_68 : _GEN_746; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_748 = 8'h45 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_69 : _GEN_747; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_749 = 8'h46 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_70 : _GEN_748; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_750 = 8'h47 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_71 : _GEN_749; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_751 = 8'h48 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_72 : _GEN_750; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_752 = 8'h49 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_73 : _GEN_751; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_753 = 8'h4a == input_0_io_dataOut_bits_0 ? io_inputs_lengths_74 : _GEN_752; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_754 = 8'h4b == input_0_io_dataOut_bits_0 ? io_inputs_lengths_75 : _GEN_753; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_755 = 8'h4c == input_0_io_dataOut_bits_0 ? io_inputs_lengths_76 : _GEN_754; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_756 = 8'h4d == input_0_io_dataOut_bits_0 ? io_inputs_lengths_77 : _GEN_755; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_757 = 8'h4e == input_0_io_dataOut_bits_0 ? io_inputs_lengths_78 : _GEN_756; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_758 = 8'h4f == input_0_io_dataOut_bits_0 ? io_inputs_lengths_79 : _GEN_757; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_759 = 8'h50 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_80 : _GEN_758; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_760 = 8'h51 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_81 : _GEN_759; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_761 = 8'h52 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_82 : _GEN_760; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_762 = 8'h53 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_83 : _GEN_761; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_763 = 8'h54 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_84 : _GEN_762; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_764 = 8'h55 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_85 : _GEN_763; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_765 = 8'h56 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_86 : _GEN_764; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_766 = 8'h57 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_87 : _GEN_765; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_767 = 8'h58 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_88 : _GEN_766; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_768 = 8'h59 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_89 : _GEN_767; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_769 = 8'h5a == input_0_io_dataOut_bits_0 ? io_inputs_lengths_90 : _GEN_768; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_770 = 8'h5b == input_0_io_dataOut_bits_0 ? io_inputs_lengths_91 : _GEN_769; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_771 = 8'h5c == input_0_io_dataOut_bits_0 ? io_inputs_lengths_92 : _GEN_770; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_772 = 8'h5d == input_0_io_dataOut_bits_0 ? io_inputs_lengths_93 : _GEN_771; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_773 = 8'h5e == input_0_io_dataOut_bits_0 ? io_inputs_lengths_94 : _GEN_772; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_774 = 8'h5f == input_0_io_dataOut_bits_0 ? io_inputs_lengths_95 : _GEN_773; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_775 = 8'h60 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_96 : _GEN_774; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_776 = 8'h61 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_97 : _GEN_775; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_777 = 8'h62 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_98 : _GEN_776; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_778 = 8'h63 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_99 : _GEN_777; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_779 = 8'h64 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_100 : _GEN_778; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_780 = 8'h65 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_101 : _GEN_779; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_781 = 8'h66 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_102 : _GEN_780; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_782 = 8'h67 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_103 : _GEN_781; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_783 = 8'h68 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_104 : _GEN_782; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_784 = 8'h69 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_105 : _GEN_783; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_785 = 8'h6a == input_0_io_dataOut_bits_0 ? io_inputs_lengths_106 : _GEN_784; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_786 = 8'h6b == input_0_io_dataOut_bits_0 ? io_inputs_lengths_107 : _GEN_785; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_787 = 8'h6c == input_0_io_dataOut_bits_0 ? io_inputs_lengths_108 : _GEN_786; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_788 = 8'h6d == input_0_io_dataOut_bits_0 ? io_inputs_lengths_109 : _GEN_787; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_789 = 8'h6e == input_0_io_dataOut_bits_0 ? io_inputs_lengths_110 : _GEN_788; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_790 = 8'h6f == input_0_io_dataOut_bits_0 ? io_inputs_lengths_111 : _GEN_789; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_791 = 8'h70 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_112 : _GEN_790; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_792 = 8'h71 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_113 : _GEN_791; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_793 = 8'h72 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_114 : _GEN_792; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_794 = 8'h73 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_115 : _GEN_793; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_795 = 8'h74 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_116 : _GEN_794; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_796 = 8'h75 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_117 : _GEN_795; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_797 = 8'h76 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_118 : _GEN_796; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_798 = 8'h77 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_119 : _GEN_797; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_799 = 8'h78 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_120 : _GEN_798; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_800 = 8'h79 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_121 : _GEN_799; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_801 = 8'h7a == input_0_io_dataOut_bits_0 ? io_inputs_lengths_122 : _GEN_800; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_802 = 8'h7b == input_0_io_dataOut_bits_0 ? io_inputs_lengths_123 : _GEN_801; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_803 = 8'h7c == input_0_io_dataOut_bits_0 ? io_inputs_lengths_124 : _GEN_802; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_804 = 8'h7d == input_0_io_dataOut_bits_0 ? io_inputs_lengths_125 : _GEN_803; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_805 = 8'h7e == input_0_io_dataOut_bits_0 ? io_inputs_lengths_126 : _GEN_804; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_806 = 8'h7f == input_0_io_dataOut_bits_0 ? io_inputs_lengths_127 : _GEN_805; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_807 = 8'h80 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_128 : _GEN_806; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_808 = 8'h81 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_129 : _GEN_807; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_809 = 8'h82 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_130 : _GEN_808; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_810 = 8'h83 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_131 : _GEN_809; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_811 = 8'h84 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_132 : _GEN_810; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_812 = 8'h85 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_133 : _GEN_811; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_813 = 8'h86 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_134 : _GEN_812; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_814 = 8'h87 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_135 : _GEN_813; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_815 = 8'h88 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_136 : _GEN_814; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_816 = 8'h89 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_137 : _GEN_815; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_817 = 8'h8a == input_0_io_dataOut_bits_0 ? io_inputs_lengths_138 : _GEN_816; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_818 = 8'h8b == input_0_io_dataOut_bits_0 ? io_inputs_lengths_139 : _GEN_817; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_819 = 8'h8c == input_0_io_dataOut_bits_0 ? io_inputs_lengths_140 : _GEN_818; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_820 = 8'h8d == input_0_io_dataOut_bits_0 ? io_inputs_lengths_141 : _GEN_819; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_821 = 8'h8e == input_0_io_dataOut_bits_0 ? io_inputs_lengths_142 : _GEN_820; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_822 = 8'h8f == input_0_io_dataOut_bits_0 ? io_inputs_lengths_143 : _GEN_821; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_823 = 8'h90 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_144 : _GEN_822; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_824 = 8'h91 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_145 : _GEN_823; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_825 = 8'h92 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_146 : _GEN_824; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_826 = 8'h93 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_147 : _GEN_825; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_827 = 8'h94 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_148 : _GEN_826; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_828 = 8'h95 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_149 : _GEN_827; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_829 = 8'h96 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_150 : _GEN_828; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_830 = 8'h97 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_151 : _GEN_829; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_831 = 8'h98 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_152 : _GEN_830; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_832 = 8'h99 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_153 : _GEN_831; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_833 = 8'h9a == input_0_io_dataOut_bits_0 ? io_inputs_lengths_154 : _GEN_832; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_834 = 8'h9b == input_0_io_dataOut_bits_0 ? io_inputs_lengths_155 : _GEN_833; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_835 = 8'h9c == input_0_io_dataOut_bits_0 ? io_inputs_lengths_156 : _GEN_834; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_836 = 8'h9d == input_0_io_dataOut_bits_0 ? io_inputs_lengths_157 : _GEN_835; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_837 = 8'h9e == input_0_io_dataOut_bits_0 ? io_inputs_lengths_158 : _GEN_836; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_838 = 8'h9f == input_0_io_dataOut_bits_0 ? io_inputs_lengths_159 : _GEN_837; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_839 = 8'ha0 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_160 : _GEN_838; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_840 = 8'ha1 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_161 : _GEN_839; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_841 = 8'ha2 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_162 : _GEN_840; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_842 = 8'ha3 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_163 : _GEN_841; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_843 = 8'ha4 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_164 : _GEN_842; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_844 = 8'ha5 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_165 : _GEN_843; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_845 = 8'ha6 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_166 : _GEN_844; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_846 = 8'ha7 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_167 : _GEN_845; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_847 = 8'ha8 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_168 : _GEN_846; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_848 = 8'ha9 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_169 : _GEN_847; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_849 = 8'haa == input_0_io_dataOut_bits_0 ? io_inputs_lengths_170 : _GEN_848; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_850 = 8'hab == input_0_io_dataOut_bits_0 ? io_inputs_lengths_171 : _GEN_849; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_851 = 8'hac == input_0_io_dataOut_bits_0 ? io_inputs_lengths_172 : _GEN_850; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_852 = 8'had == input_0_io_dataOut_bits_0 ? io_inputs_lengths_173 : _GEN_851; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_853 = 8'hae == input_0_io_dataOut_bits_0 ? io_inputs_lengths_174 : _GEN_852; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_854 = 8'haf == input_0_io_dataOut_bits_0 ? io_inputs_lengths_175 : _GEN_853; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_855 = 8'hb0 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_176 : _GEN_854; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_856 = 8'hb1 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_177 : _GEN_855; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_857 = 8'hb2 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_178 : _GEN_856; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_858 = 8'hb3 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_179 : _GEN_857; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_859 = 8'hb4 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_180 : _GEN_858; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_860 = 8'hb5 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_181 : _GEN_859; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_861 = 8'hb6 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_182 : _GEN_860; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_862 = 8'hb7 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_183 : _GEN_861; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_863 = 8'hb8 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_184 : _GEN_862; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_864 = 8'hb9 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_185 : _GEN_863; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_865 = 8'hba == input_0_io_dataOut_bits_0 ? io_inputs_lengths_186 : _GEN_864; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_866 = 8'hbb == input_0_io_dataOut_bits_0 ? io_inputs_lengths_187 : _GEN_865; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_867 = 8'hbc == input_0_io_dataOut_bits_0 ? io_inputs_lengths_188 : _GEN_866; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_868 = 8'hbd == input_0_io_dataOut_bits_0 ? io_inputs_lengths_189 : _GEN_867; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_869 = 8'hbe == input_0_io_dataOut_bits_0 ? io_inputs_lengths_190 : _GEN_868; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_870 = 8'hbf == input_0_io_dataOut_bits_0 ? io_inputs_lengths_191 : _GEN_869; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_871 = 8'hc0 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_192 : _GEN_870; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_872 = 8'hc1 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_193 : _GEN_871; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_873 = 8'hc2 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_194 : _GEN_872; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_874 = 8'hc3 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_195 : _GEN_873; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_875 = 8'hc4 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_196 : _GEN_874; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_876 = 8'hc5 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_197 : _GEN_875; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_877 = 8'hc6 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_198 : _GEN_876; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_878 = 8'hc7 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_199 : _GEN_877; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_879 = 8'hc8 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_200 : _GEN_878; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_880 = 8'hc9 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_201 : _GEN_879; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_881 = 8'hca == input_0_io_dataOut_bits_0 ? io_inputs_lengths_202 : _GEN_880; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_882 = 8'hcb == input_0_io_dataOut_bits_0 ? io_inputs_lengths_203 : _GEN_881; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_883 = 8'hcc == input_0_io_dataOut_bits_0 ? io_inputs_lengths_204 : _GEN_882; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_884 = 8'hcd == input_0_io_dataOut_bits_0 ? io_inputs_lengths_205 : _GEN_883; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_885 = 8'hce == input_0_io_dataOut_bits_0 ? io_inputs_lengths_206 : _GEN_884; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_886 = 8'hcf == input_0_io_dataOut_bits_0 ? io_inputs_lengths_207 : _GEN_885; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_887 = 8'hd0 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_208 : _GEN_886; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_888 = 8'hd1 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_209 : _GEN_887; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_889 = 8'hd2 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_210 : _GEN_888; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_890 = 8'hd3 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_211 : _GEN_889; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_891 = 8'hd4 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_212 : _GEN_890; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_892 = 8'hd5 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_213 : _GEN_891; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_893 = 8'hd6 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_214 : _GEN_892; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_894 = 8'hd7 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_215 : _GEN_893; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_895 = 8'hd8 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_216 : _GEN_894; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_896 = 8'hd9 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_217 : _GEN_895; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_897 = 8'hda == input_0_io_dataOut_bits_0 ? io_inputs_lengths_218 : _GEN_896; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_898 = 8'hdb == input_0_io_dataOut_bits_0 ? io_inputs_lengths_219 : _GEN_897; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_899 = 8'hdc == input_0_io_dataOut_bits_0 ? io_inputs_lengths_220 : _GEN_898; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_900 = 8'hdd == input_0_io_dataOut_bits_0 ? io_inputs_lengths_221 : _GEN_899; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_901 = 8'hde == input_0_io_dataOut_bits_0 ? io_inputs_lengths_222 : _GEN_900; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_902 = 8'hdf == input_0_io_dataOut_bits_0 ? io_inputs_lengths_223 : _GEN_901; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_903 = 8'he0 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_224 : _GEN_902; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_904 = 8'he1 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_225 : _GEN_903; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_905 = 8'he2 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_226 : _GEN_904; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_906 = 8'he3 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_227 : _GEN_905; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_907 = 8'he4 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_228 : _GEN_906; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_908 = 8'he5 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_229 : _GEN_907; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_909 = 8'he6 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_230 : _GEN_908; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_910 = 8'he7 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_231 : _GEN_909; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_911 = 8'he8 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_232 : _GEN_910; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_912 = 8'he9 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_233 : _GEN_911; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_913 = 8'hea == input_0_io_dataOut_bits_0 ? io_inputs_lengths_234 : _GEN_912; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_914 = 8'heb == input_0_io_dataOut_bits_0 ? io_inputs_lengths_235 : _GEN_913; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_915 = 8'hec == input_0_io_dataOut_bits_0 ? io_inputs_lengths_236 : _GEN_914; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_916 = 8'hed == input_0_io_dataOut_bits_0 ? io_inputs_lengths_237 : _GEN_915; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_917 = 8'hee == input_0_io_dataOut_bits_0 ? io_inputs_lengths_238 : _GEN_916; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_918 = 8'hef == input_0_io_dataOut_bits_0 ? io_inputs_lengths_239 : _GEN_917; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_919 = 8'hf0 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_240 : _GEN_918; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_920 = 8'hf1 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_241 : _GEN_919; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_921 = 8'hf2 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_242 : _GEN_920; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_922 = 8'hf3 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_243 : _GEN_921; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_923 = 8'hf4 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_244 : _GEN_922; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_924 = 8'hf5 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_245 : _GEN_923; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_925 = 8'hf6 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_246 : _GEN_924; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_926 = 8'hf7 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_247 : _GEN_925; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_927 = 8'hf8 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_248 : _GEN_926; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_928 = 8'hf9 == input_0_io_dataOut_bits_0 ? io_inputs_lengths_249 : _GEN_927; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_929 = 8'hfa == input_0_io_dataOut_bits_0 ? io_inputs_lengths_250 : _GEN_928; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_930 = 8'hfb == input_0_io_dataOut_bits_0 ? io_inputs_lengths_251 : _GEN_929; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_931 = 8'hfc == input_0_io_dataOut_bits_0 ? io_inputs_lengths_252 : _GEN_930; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_932 = 8'hfd == input_0_io_dataOut_bits_0 ? io_inputs_lengths_253 : _GEN_931; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_933 = 8'hfe == input_0_io_dataOut_bits_0 ? io_inputs_lengths_254 : _GEN_932; // @[compressorOutput.scala 143:42]
  wire [4:0] _GEN_934 = 8'hff == input_0_io_dataOut_bits_0 ? io_inputs_lengths_255 : _GEN_933; // @[compressorOutput.scala 143:42]
  wire [4:0] _T_30 = 5'h1c - _GEN_934; // @[compressorOutput.scala 145:95]
  wire [23:0] _GEN_936 = 8'h1 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_1 : io_inputs_codewords_0; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_937 = 8'h2 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_2 : _GEN_936; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_938 = 8'h3 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_3 : _GEN_937; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_939 = 8'h4 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_4 : _GEN_938; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_940 = 8'h5 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_5 : _GEN_939; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_941 = 8'h6 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_6 : _GEN_940; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_942 = 8'h7 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_7 : _GEN_941; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_943 = 8'h8 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_8 : _GEN_942; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_944 = 8'h9 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_9 : _GEN_943; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_945 = 8'ha == input_0_io_dataOut_bits_0 ? io_inputs_codewords_10 : _GEN_944; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_946 = 8'hb == input_0_io_dataOut_bits_0 ? io_inputs_codewords_11 : _GEN_945; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_947 = 8'hc == input_0_io_dataOut_bits_0 ? io_inputs_codewords_12 : _GEN_946; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_948 = 8'hd == input_0_io_dataOut_bits_0 ? io_inputs_codewords_13 : _GEN_947; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_949 = 8'he == input_0_io_dataOut_bits_0 ? io_inputs_codewords_14 : _GEN_948; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_950 = 8'hf == input_0_io_dataOut_bits_0 ? io_inputs_codewords_15 : _GEN_949; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_951 = 8'h10 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_16 : _GEN_950; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_952 = 8'h11 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_17 : _GEN_951; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_953 = 8'h12 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_18 : _GEN_952; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_954 = 8'h13 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_19 : _GEN_953; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_955 = 8'h14 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_20 : _GEN_954; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_956 = 8'h15 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_21 : _GEN_955; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_957 = 8'h16 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_22 : _GEN_956; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_958 = 8'h17 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_23 : _GEN_957; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_959 = 8'h18 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_24 : _GEN_958; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_960 = 8'h19 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_25 : _GEN_959; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_961 = 8'h1a == input_0_io_dataOut_bits_0 ? io_inputs_codewords_26 : _GEN_960; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_962 = 8'h1b == input_0_io_dataOut_bits_0 ? io_inputs_codewords_27 : _GEN_961; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_963 = 8'h1c == input_0_io_dataOut_bits_0 ? io_inputs_codewords_28 : _GEN_962; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_964 = 8'h1d == input_0_io_dataOut_bits_0 ? io_inputs_codewords_29 : _GEN_963; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_965 = 8'h1e == input_0_io_dataOut_bits_0 ? io_inputs_codewords_30 : _GEN_964; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_966 = 8'h1f == input_0_io_dataOut_bits_0 ? io_inputs_codewords_31 : _GEN_965; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_967 = 8'h20 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_32 : _GEN_966; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_968 = 8'h21 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_33 : _GEN_967; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_969 = 8'h22 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_34 : _GEN_968; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_970 = 8'h23 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_35 : _GEN_969; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_971 = 8'h24 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_36 : _GEN_970; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_972 = 8'h25 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_37 : _GEN_971; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_973 = 8'h26 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_38 : _GEN_972; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_974 = 8'h27 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_39 : _GEN_973; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_975 = 8'h28 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_40 : _GEN_974; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_976 = 8'h29 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_41 : _GEN_975; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_977 = 8'h2a == input_0_io_dataOut_bits_0 ? io_inputs_codewords_42 : _GEN_976; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_978 = 8'h2b == input_0_io_dataOut_bits_0 ? io_inputs_codewords_43 : _GEN_977; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_979 = 8'h2c == input_0_io_dataOut_bits_0 ? io_inputs_codewords_44 : _GEN_978; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_980 = 8'h2d == input_0_io_dataOut_bits_0 ? io_inputs_codewords_45 : _GEN_979; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_981 = 8'h2e == input_0_io_dataOut_bits_0 ? io_inputs_codewords_46 : _GEN_980; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_982 = 8'h2f == input_0_io_dataOut_bits_0 ? io_inputs_codewords_47 : _GEN_981; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_983 = 8'h30 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_48 : _GEN_982; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_984 = 8'h31 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_49 : _GEN_983; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_985 = 8'h32 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_50 : _GEN_984; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_986 = 8'h33 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_51 : _GEN_985; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_987 = 8'h34 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_52 : _GEN_986; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_988 = 8'h35 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_53 : _GEN_987; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_989 = 8'h36 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_54 : _GEN_988; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_990 = 8'h37 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_55 : _GEN_989; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_991 = 8'h38 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_56 : _GEN_990; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_992 = 8'h39 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_57 : _GEN_991; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_993 = 8'h3a == input_0_io_dataOut_bits_0 ? io_inputs_codewords_58 : _GEN_992; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_994 = 8'h3b == input_0_io_dataOut_bits_0 ? io_inputs_codewords_59 : _GEN_993; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_995 = 8'h3c == input_0_io_dataOut_bits_0 ? io_inputs_codewords_60 : _GEN_994; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_996 = 8'h3d == input_0_io_dataOut_bits_0 ? io_inputs_codewords_61 : _GEN_995; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_997 = 8'h3e == input_0_io_dataOut_bits_0 ? io_inputs_codewords_62 : _GEN_996; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_998 = 8'h3f == input_0_io_dataOut_bits_0 ? io_inputs_codewords_63 : _GEN_997; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_999 = 8'h40 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_64 : _GEN_998; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1000 = 8'h41 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_65 : _GEN_999; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1001 = 8'h42 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_66 : _GEN_1000; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1002 = 8'h43 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_67 : _GEN_1001; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1003 = 8'h44 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_68 : _GEN_1002; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1004 = 8'h45 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_69 : _GEN_1003; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1005 = 8'h46 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_70 : _GEN_1004; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1006 = 8'h47 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_71 : _GEN_1005; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1007 = 8'h48 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_72 : _GEN_1006; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1008 = 8'h49 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_73 : _GEN_1007; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1009 = 8'h4a == input_0_io_dataOut_bits_0 ? io_inputs_codewords_74 : _GEN_1008; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1010 = 8'h4b == input_0_io_dataOut_bits_0 ? io_inputs_codewords_75 : _GEN_1009; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1011 = 8'h4c == input_0_io_dataOut_bits_0 ? io_inputs_codewords_76 : _GEN_1010; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1012 = 8'h4d == input_0_io_dataOut_bits_0 ? io_inputs_codewords_77 : _GEN_1011; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1013 = 8'h4e == input_0_io_dataOut_bits_0 ? io_inputs_codewords_78 : _GEN_1012; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1014 = 8'h4f == input_0_io_dataOut_bits_0 ? io_inputs_codewords_79 : _GEN_1013; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1015 = 8'h50 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_80 : _GEN_1014; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1016 = 8'h51 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_81 : _GEN_1015; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1017 = 8'h52 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_82 : _GEN_1016; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1018 = 8'h53 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_83 : _GEN_1017; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1019 = 8'h54 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_84 : _GEN_1018; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1020 = 8'h55 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_85 : _GEN_1019; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1021 = 8'h56 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_86 : _GEN_1020; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1022 = 8'h57 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_87 : _GEN_1021; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1023 = 8'h58 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_88 : _GEN_1022; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1024 = 8'h59 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_89 : _GEN_1023; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1025 = 8'h5a == input_0_io_dataOut_bits_0 ? io_inputs_codewords_90 : _GEN_1024; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1026 = 8'h5b == input_0_io_dataOut_bits_0 ? io_inputs_codewords_91 : _GEN_1025; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1027 = 8'h5c == input_0_io_dataOut_bits_0 ? io_inputs_codewords_92 : _GEN_1026; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1028 = 8'h5d == input_0_io_dataOut_bits_0 ? io_inputs_codewords_93 : _GEN_1027; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1029 = 8'h5e == input_0_io_dataOut_bits_0 ? io_inputs_codewords_94 : _GEN_1028; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1030 = 8'h5f == input_0_io_dataOut_bits_0 ? io_inputs_codewords_95 : _GEN_1029; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1031 = 8'h60 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_96 : _GEN_1030; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1032 = 8'h61 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_97 : _GEN_1031; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1033 = 8'h62 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_98 : _GEN_1032; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1034 = 8'h63 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_99 : _GEN_1033; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1035 = 8'h64 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_100 : _GEN_1034; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1036 = 8'h65 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_101 : _GEN_1035; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1037 = 8'h66 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_102 : _GEN_1036; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1038 = 8'h67 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_103 : _GEN_1037; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1039 = 8'h68 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_104 : _GEN_1038; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1040 = 8'h69 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_105 : _GEN_1039; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1041 = 8'h6a == input_0_io_dataOut_bits_0 ? io_inputs_codewords_106 : _GEN_1040; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1042 = 8'h6b == input_0_io_dataOut_bits_0 ? io_inputs_codewords_107 : _GEN_1041; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1043 = 8'h6c == input_0_io_dataOut_bits_0 ? io_inputs_codewords_108 : _GEN_1042; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1044 = 8'h6d == input_0_io_dataOut_bits_0 ? io_inputs_codewords_109 : _GEN_1043; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1045 = 8'h6e == input_0_io_dataOut_bits_0 ? io_inputs_codewords_110 : _GEN_1044; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1046 = 8'h6f == input_0_io_dataOut_bits_0 ? io_inputs_codewords_111 : _GEN_1045; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1047 = 8'h70 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_112 : _GEN_1046; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1048 = 8'h71 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_113 : _GEN_1047; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1049 = 8'h72 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_114 : _GEN_1048; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1050 = 8'h73 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_115 : _GEN_1049; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1051 = 8'h74 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_116 : _GEN_1050; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1052 = 8'h75 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_117 : _GEN_1051; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1053 = 8'h76 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_118 : _GEN_1052; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1054 = 8'h77 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_119 : _GEN_1053; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1055 = 8'h78 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_120 : _GEN_1054; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1056 = 8'h79 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_121 : _GEN_1055; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1057 = 8'h7a == input_0_io_dataOut_bits_0 ? io_inputs_codewords_122 : _GEN_1056; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1058 = 8'h7b == input_0_io_dataOut_bits_0 ? io_inputs_codewords_123 : _GEN_1057; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1059 = 8'h7c == input_0_io_dataOut_bits_0 ? io_inputs_codewords_124 : _GEN_1058; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1060 = 8'h7d == input_0_io_dataOut_bits_0 ? io_inputs_codewords_125 : _GEN_1059; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1061 = 8'h7e == input_0_io_dataOut_bits_0 ? io_inputs_codewords_126 : _GEN_1060; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1062 = 8'h7f == input_0_io_dataOut_bits_0 ? io_inputs_codewords_127 : _GEN_1061; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1063 = 8'h80 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_128 : _GEN_1062; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1064 = 8'h81 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_129 : _GEN_1063; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1065 = 8'h82 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_130 : _GEN_1064; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1066 = 8'h83 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_131 : _GEN_1065; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1067 = 8'h84 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_132 : _GEN_1066; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1068 = 8'h85 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_133 : _GEN_1067; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1069 = 8'h86 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_134 : _GEN_1068; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1070 = 8'h87 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_135 : _GEN_1069; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1071 = 8'h88 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_136 : _GEN_1070; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1072 = 8'h89 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_137 : _GEN_1071; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1073 = 8'h8a == input_0_io_dataOut_bits_0 ? io_inputs_codewords_138 : _GEN_1072; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1074 = 8'h8b == input_0_io_dataOut_bits_0 ? io_inputs_codewords_139 : _GEN_1073; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1075 = 8'h8c == input_0_io_dataOut_bits_0 ? io_inputs_codewords_140 : _GEN_1074; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1076 = 8'h8d == input_0_io_dataOut_bits_0 ? io_inputs_codewords_141 : _GEN_1075; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1077 = 8'h8e == input_0_io_dataOut_bits_0 ? io_inputs_codewords_142 : _GEN_1076; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1078 = 8'h8f == input_0_io_dataOut_bits_0 ? io_inputs_codewords_143 : _GEN_1077; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1079 = 8'h90 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_144 : _GEN_1078; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1080 = 8'h91 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_145 : _GEN_1079; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1081 = 8'h92 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_146 : _GEN_1080; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1082 = 8'h93 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_147 : _GEN_1081; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1083 = 8'h94 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_148 : _GEN_1082; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1084 = 8'h95 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_149 : _GEN_1083; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1085 = 8'h96 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_150 : _GEN_1084; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1086 = 8'h97 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_151 : _GEN_1085; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1087 = 8'h98 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_152 : _GEN_1086; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1088 = 8'h99 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_153 : _GEN_1087; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1089 = 8'h9a == input_0_io_dataOut_bits_0 ? io_inputs_codewords_154 : _GEN_1088; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1090 = 8'h9b == input_0_io_dataOut_bits_0 ? io_inputs_codewords_155 : _GEN_1089; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1091 = 8'h9c == input_0_io_dataOut_bits_0 ? io_inputs_codewords_156 : _GEN_1090; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1092 = 8'h9d == input_0_io_dataOut_bits_0 ? io_inputs_codewords_157 : _GEN_1091; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1093 = 8'h9e == input_0_io_dataOut_bits_0 ? io_inputs_codewords_158 : _GEN_1092; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1094 = 8'h9f == input_0_io_dataOut_bits_0 ? io_inputs_codewords_159 : _GEN_1093; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1095 = 8'ha0 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_160 : _GEN_1094; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1096 = 8'ha1 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_161 : _GEN_1095; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1097 = 8'ha2 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_162 : _GEN_1096; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1098 = 8'ha3 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_163 : _GEN_1097; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1099 = 8'ha4 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_164 : _GEN_1098; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1100 = 8'ha5 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_165 : _GEN_1099; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1101 = 8'ha6 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_166 : _GEN_1100; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1102 = 8'ha7 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_167 : _GEN_1101; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1103 = 8'ha8 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_168 : _GEN_1102; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1104 = 8'ha9 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_169 : _GEN_1103; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1105 = 8'haa == input_0_io_dataOut_bits_0 ? io_inputs_codewords_170 : _GEN_1104; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1106 = 8'hab == input_0_io_dataOut_bits_0 ? io_inputs_codewords_171 : _GEN_1105; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1107 = 8'hac == input_0_io_dataOut_bits_0 ? io_inputs_codewords_172 : _GEN_1106; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1108 = 8'had == input_0_io_dataOut_bits_0 ? io_inputs_codewords_173 : _GEN_1107; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1109 = 8'hae == input_0_io_dataOut_bits_0 ? io_inputs_codewords_174 : _GEN_1108; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1110 = 8'haf == input_0_io_dataOut_bits_0 ? io_inputs_codewords_175 : _GEN_1109; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1111 = 8'hb0 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_176 : _GEN_1110; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1112 = 8'hb1 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_177 : _GEN_1111; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1113 = 8'hb2 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_178 : _GEN_1112; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1114 = 8'hb3 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_179 : _GEN_1113; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1115 = 8'hb4 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_180 : _GEN_1114; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1116 = 8'hb5 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_181 : _GEN_1115; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1117 = 8'hb6 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_182 : _GEN_1116; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1118 = 8'hb7 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_183 : _GEN_1117; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1119 = 8'hb8 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_184 : _GEN_1118; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1120 = 8'hb9 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_185 : _GEN_1119; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1121 = 8'hba == input_0_io_dataOut_bits_0 ? io_inputs_codewords_186 : _GEN_1120; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1122 = 8'hbb == input_0_io_dataOut_bits_0 ? io_inputs_codewords_187 : _GEN_1121; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1123 = 8'hbc == input_0_io_dataOut_bits_0 ? io_inputs_codewords_188 : _GEN_1122; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1124 = 8'hbd == input_0_io_dataOut_bits_0 ? io_inputs_codewords_189 : _GEN_1123; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1125 = 8'hbe == input_0_io_dataOut_bits_0 ? io_inputs_codewords_190 : _GEN_1124; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1126 = 8'hbf == input_0_io_dataOut_bits_0 ? io_inputs_codewords_191 : _GEN_1125; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1127 = 8'hc0 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_192 : _GEN_1126; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1128 = 8'hc1 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_193 : _GEN_1127; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1129 = 8'hc2 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_194 : _GEN_1128; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1130 = 8'hc3 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_195 : _GEN_1129; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1131 = 8'hc4 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_196 : _GEN_1130; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1132 = 8'hc5 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_197 : _GEN_1131; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1133 = 8'hc6 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_198 : _GEN_1132; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1134 = 8'hc7 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_199 : _GEN_1133; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1135 = 8'hc8 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_200 : _GEN_1134; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1136 = 8'hc9 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_201 : _GEN_1135; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1137 = 8'hca == input_0_io_dataOut_bits_0 ? io_inputs_codewords_202 : _GEN_1136; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1138 = 8'hcb == input_0_io_dataOut_bits_0 ? io_inputs_codewords_203 : _GEN_1137; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1139 = 8'hcc == input_0_io_dataOut_bits_0 ? io_inputs_codewords_204 : _GEN_1138; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1140 = 8'hcd == input_0_io_dataOut_bits_0 ? io_inputs_codewords_205 : _GEN_1139; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1141 = 8'hce == input_0_io_dataOut_bits_0 ? io_inputs_codewords_206 : _GEN_1140; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1142 = 8'hcf == input_0_io_dataOut_bits_0 ? io_inputs_codewords_207 : _GEN_1141; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1143 = 8'hd0 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_208 : _GEN_1142; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1144 = 8'hd1 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_209 : _GEN_1143; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1145 = 8'hd2 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_210 : _GEN_1144; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1146 = 8'hd3 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_211 : _GEN_1145; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1147 = 8'hd4 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_212 : _GEN_1146; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1148 = 8'hd5 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_213 : _GEN_1147; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1149 = 8'hd6 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_214 : _GEN_1148; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1150 = 8'hd7 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_215 : _GEN_1149; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1151 = 8'hd8 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_216 : _GEN_1150; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1152 = 8'hd9 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_217 : _GEN_1151; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1153 = 8'hda == input_0_io_dataOut_bits_0 ? io_inputs_codewords_218 : _GEN_1152; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1154 = 8'hdb == input_0_io_dataOut_bits_0 ? io_inputs_codewords_219 : _GEN_1153; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1155 = 8'hdc == input_0_io_dataOut_bits_0 ? io_inputs_codewords_220 : _GEN_1154; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1156 = 8'hdd == input_0_io_dataOut_bits_0 ? io_inputs_codewords_221 : _GEN_1155; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1157 = 8'hde == input_0_io_dataOut_bits_0 ? io_inputs_codewords_222 : _GEN_1156; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1158 = 8'hdf == input_0_io_dataOut_bits_0 ? io_inputs_codewords_223 : _GEN_1157; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1159 = 8'he0 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_224 : _GEN_1158; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1160 = 8'he1 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_225 : _GEN_1159; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1161 = 8'he2 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_226 : _GEN_1160; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1162 = 8'he3 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_227 : _GEN_1161; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1163 = 8'he4 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_228 : _GEN_1162; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1164 = 8'he5 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_229 : _GEN_1163; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1165 = 8'he6 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_230 : _GEN_1164; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1166 = 8'he7 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_231 : _GEN_1165; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1167 = 8'he8 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_232 : _GEN_1166; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1168 = 8'he9 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_233 : _GEN_1167; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1169 = 8'hea == input_0_io_dataOut_bits_0 ? io_inputs_codewords_234 : _GEN_1168; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1170 = 8'heb == input_0_io_dataOut_bits_0 ? io_inputs_codewords_235 : _GEN_1169; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1171 = 8'hec == input_0_io_dataOut_bits_0 ? io_inputs_codewords_236 : _GEN_1170; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1172 = 8'hed == input_0_io_dataOut_bits_0 ? io_inputs_codewords_237 : _GEN_1171; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1173 = 8'hee == input_0_io_dataOut_bits_0 ? io_inputs_codewords_238 : _GEN_1172; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1174 = 8'hef == input_0_io_dataOut_bits_0 ? io_inputs_codewords_239 : _GEN_1173; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1175 = 8'hf0 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_240 : _GEN_1174; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1176 = 8'hf1 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_241 : _GEN_1175; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1177 = 8'hf2 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_242 : _GEN_1176; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1178 = 8'hf3 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_243 : _GEN_1177; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1179 = 8'hf4 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_244 : _GEN_1178; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1180 = 8'hf5 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_245 : _GEN_1179; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1181 = 8'hf6 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_246 : _GEN_1180; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1182 = 8'hf7 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_247 : _GEN_1181; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1183 = 8'hf8 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_248 : _GEN_1182; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1184 = 8'hf9 == input_0_io_dataOut_bits_0 ? io_inputs_codewords_249 : _GEN_1183; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1185 = 8'hfa == input_0_io_dataOut_bits_0 ? io_inputs_codewords_250 : _GEN_1184; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1186 = 8'hfb == input_0_io_dataOut_bits_0 ? io_inputs_codewords_251 : _GEN_1185; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1187 = 8'hfc == input_0_io_dataOut_bits_0 ? io_inputs_codewords_252 : _GEN_1186; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1188 = 8'hfd == input_0_io_dataOut_bits_0 ? io_inputs_codewords_253 : _GEN_1187; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1189 = 8'hfe == input_0_io_dataOut_bits_0 ? io_inputs_codewords_254 : _GEN_1188; // @[compressorOutput.scala 145:59]
  wire [23:0] _GEN_1190 = 8'hff == input_0_io_dataOut_bits_0 ? io_inputs_codewords_255 : _GEN_1189; // @[compressorOutput.scala 145:59]
  wire [54:0] _GEN_1223 = {{31'd0}, _GEN_1190}; // @[compressorOutput.scala 145:59]
  wire [54:0] _T_31 = _GEN_1223 << _T_30; // @[compressorOutput.scala 145:59]
  wire  _GEN_1192 = input_0_io_dataOut_valid; // @[compressorOutput.scala 141:47]
  wire [4:0] _GEN_1193 = input_0_io_dataOut_valid ? _GEN_934 : 5'h0; // @[compressorOutput.scala 141:47]
  wire [54:0] _GEN_1194 = input_0_io_dataOut_valid ? _T_31 : 55'h0; // @[compressorOutput.scala 141:47]
  wire  _GEN_1196 = _T_25 & _GEN_1192; // @[compressorOutput.scala 140:63]
  wire [4:0] _GEN_1197 = _T_25 ? _GEN_1193 : 5'h0; // @[compressorOutput.scala 140:63]
  wire [54:0] _GEN_1198 = _T_25 ? _GEN_1194 : 55'h0; // @[compressorOutput.scala 140:63]
  wire  _T_34 = iterations_0 >= 13'h1000; // @[compressorOutput.scala 158:29]
  wire  _GEN_1201 = _T_24 & _T_25; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_1202 = _T_24 ? _T_26[12:0] : 13'h0; // @[Conditional.scala 39:67]
  wire  _GEN_1203 = _T_24 & _GEN_1196; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_1204 = _T_24 ? _GEN_1197 : 5'h0; // @[Conditional.scala 39:67]
  wire [54:0] _GEN_1205 = _T_24 ? _GEN_1198 : 55'h0; // @[Conditional.scala 39:67]
  wire  _GEN_1208 = _T_1 ? 1'h0 : _GEN_1201; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_1209 = _T_1 ? 13'h0 : _GEN_1202; // @[Conditional.scala 39:67]
  wire  _GEN_1210 = _T_1 | _GEN_1203; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_1211 = _T_1 ? 5'h1c : _GEN_1204; // @[Conditional.scala 39:67]
  wire [54:0] _GEN_1212 = _T_1 ? {{27'd0}, _GEN_674} : _GEN_1205; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_1218 = _T ? 13'h0 : _GEN_1209; // @[Conditional.scala 40:58]
  wire [54:0] _GEN_1221 = _T ? 55'h0 : _GEN_1212; // @[Conditional.scala 40:58]
  compressorInput input_0 ( // @[compressorOutput.scala 34:51]
    .io_input_currentByteOut(input_0_io_input_currentByteOut),
    .io_input_dataIn_0(input_0_io_input_dataIn_0),
    .io_input_valid(input_0_io_input_valid),
    .io_input_ready(input_0_io_input_ready),
    .io_currentByte(input_0_io_currentByte),
    .io_dataOut_ready(input_0_io_dataOut_ready),
    .io_dataOut_valid(input_0_io_dataOut_valid),
    .io_dataOut_bits_0(input_0_io_dataOut_bits_0)
  );
  assign io_dataIn_0_currentByteOut = input_0_io_input_currentByteOut; // @[compressorOutput.scala 54:27]
  assign io_dataIn_0_ready = input_0_io_input_ready; // @[compressorOutput.scala 54:27]
  assign io_outputs_0_dataOut = _GEN_1221[27:0]; // @[compressorOutput.scala 49:31 compressorOutput.scala 92:33 compressorOutput.scala 101:33 compressorOutput.scala 117:31 compressorOutput.scala 139:35 compressorOutput.scala 144:39]
  assign io_outputs_0_dataLength = _T ? 5'h0 : _GEN_1211; // @[compressorOutput.scala 51:34 compressorOutput.scala 85:32 compressorOutput.scala 138:38 compressorOutput.scala 143:42]
  assign io_outputs_0_valid = _T ? 1'h0 : _GEN_1210; // @[compressorOutput.scala 50:29 compressorOutput.scala 84:27 compressorOutput.scala 137:33 compressorOutput.scala 142:37]
  assign io_finished = state == 2'h0; // @[compressorOutput.scala 165:15]
  assign input_0_io_input_dataIn_0 = io_dataIn_0_dataIn_0; // @[compressorOutput.scala 54:27]
  assign input_0_io_input_valid = io_dataIn_0_valid; // @[compressorOutput.scala 54:27]
  assign input_0_io_currentByte = _GEN_1218[11:0]; // @[compressorOutput.scala 53:33 compressorOutput.scala 73:37 compressorOutput.scala 136:37]
  assign input_0_io_dataOut_ready = _T ? 1'h0 : _GEN_1208; // @[compressorOutput.scala 52:35 compressorOutput.scala 72:39 compressorOutput.scala 135:39]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  iterations_0 = _RAND_1[12:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T) begin
      if (io_start) begin
        state <= 2'h1;
      end
    end else if (_T_1) begin
      if (io_outputs_0_ready) begin
        if (_T_23) begin
          state <= 2'h2;
        end
      end
    end else if (_T_24) begin
      if (_T_34) begin
        state <= 2'h0;
      end
    end
    if (_T) begin
      iterations_0 <= 13'h0;
    end else if (_T_1) begin
      if (io_outputs_0_ready) begin
        if (_T_23) begin
          iterations_0 <= 13'h0;
        end else begin
          iterations_0 <= _T_20;
        end
      end
    end else if (_T_24) begin
      if (_T_25) begin
        if (input_0_io_dataOut_valid) begin
          if (io_outputs_0_ready) begin
            iterations_0 <= _T_20;
          end
        end
      end
    end
  end
endmodule
module topLevel(
  input         clock,
  input         reset,
  input         io_start,
  output [11:0] io_characterFrequencyInputs_currentByteOut,
  input  [7:0]  io_characterFrequencyInputs_dataIn_0,
  input         io_characterFrequencyInputs_valid,
  output        io_characterFrequencyInputs_ready,
  output [11:0] io_compressionInputs_0_currentByteOut,
  input  [7:0]  io_compressionInputs_0_dataIn_0,
  input         io_compressionInputs_0_valid,
  output        io_compressionInputs_0_ready,
  output [27:0] io_outputs_0_dataOut,
  output [4:0]  io_outputs_0_dataLength,
  output        io_outputs_0_valid,
  input         io_outputs_0_ready,
  output        io_finished
);
  wire  cfm_clock; // @[topLevel.scala 55:19]
  wire  cfm_reset; // @[topLevel.scala 55:19]
  wire  cfm_io_start; // @[topLevel.scala 55:19]
  wire [11:0] cfm_io_input_currentByteOut; // @[topLevel.scala 55:19]
  wire [7:0] cfm_io_input_dataIn_0; // @[topLevel.scala 55:19]
  wire  cfm_io_input_valid; // @[topLevel.scala 55:19]
  wire  cfm_io_input_ready; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_0; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_1; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_2; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_3; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_4; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_5; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_6; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_7; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_8; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_9; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_10; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_11; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_12; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_13; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_14; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_15; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_16; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_17; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_18; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_19; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_20; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_21; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_22; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_23; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_24; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_25; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_26; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_27; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_28; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_29; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_30; // @[topLevel.scala 55:19]
  wire [12:0] cfm_io_outputs_sortedFrequency_31; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_0; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_1; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_2; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_3; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_4; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_5; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_6; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_7; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_8; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_9; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_10; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_11; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_12; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_13; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_14; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_15; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_16; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_17; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_18; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_19; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_20; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_21; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_22; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_23; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_24; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_25; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_26; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_27; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_28; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_29; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_30; // @[topLevel.scala 55:19]
  wire [8:0] cfm_io_outputs_sortedCharacter_31; // @[topLevel.scala 55:19]
  wire  cfm_io_finished; // @[topLevel.scala 55:19]
  wire  tg_clock; // @[topLevel.scala 56:18]
  wire  tg_reset; // @[topLevel.scala 56:18]
  wire  tg_io_start; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_0; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_1; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_2; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_3; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_4; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_5; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_6; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_7; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_8; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_9; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_10; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_11; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_12; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_13; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_14; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_15; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_16; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_17; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_18; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_19; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_20; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_21; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_22; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_23; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_24; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_25; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_26; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_27; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_28; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_29; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_30; // @[topLevel.scala 56:18]
  wire [12:0] tg_io_inputs_sortedFrequency_31; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_0; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_1; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_2; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_3; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_4; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_5; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_6; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_7; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_8; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_9; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_10; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_11; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_12; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_13; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_14; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_15; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_16; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_17; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_18; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_19; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_20; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_21; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_22; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_23; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_24; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_25; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_26; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_27; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_28; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_29; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_30; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_inputs_sortedCharacter_31; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_0; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_1; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_2; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_3; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_4; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_5; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_6; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_7; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_8; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_9; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_10; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_11; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_12; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_13; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_14; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_15; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_16; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_17; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_18; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_19; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_20; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_21; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_22; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_23; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_24; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_25; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_26; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_27; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_28; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_29; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_30; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_31; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_32; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_33; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_34; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_35; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_36; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_37; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_38; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_39; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_40; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_41; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_42; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_43; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_44; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_45; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_46; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_47; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_48; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_49; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_50; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_51; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_52; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_53; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_54; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_55; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_56; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_57; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_58; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_59; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_60; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_61; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_62; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_leftNode_63; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_0; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_1; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_2; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_3; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_4; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_5; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_6; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_7; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_8; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_9; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_10; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_11; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_12; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_13; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_14; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_15; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_16; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_17; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_18; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_19; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_20; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_21; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_22; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_23; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_24; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_25; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_26; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_27; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_28; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_29; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_30; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_31; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_32; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_33; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_34; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_35; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_36; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_37; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_38; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_39; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_40; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_41; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_42; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_43; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_44; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_45; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_46; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_47; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_48; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_49; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_50; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_51; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_52; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_53; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_54; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_55; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_56; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_57; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_58; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_59; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_60; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_61; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_62; // @[topLevel.scala 56:18]
  wire [8:0] tg_io_outputs_rightNode_63; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_0; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_1; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_2; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_3; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_4; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_5; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_6; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_7; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_8; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_9; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_10; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_11; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_12; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_13; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_14; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_15; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_16; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_17; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_18; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_19; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_20; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_21; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_22; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_23; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_24; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_25; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_26; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_27; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_28; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_29; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_30; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_31; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_32; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_33; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_34; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_35; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_36; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_37; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_38; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_39; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_40; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_41; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_42; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_43; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_44; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_45; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_46; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_47; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_48; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_49; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_50; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_51; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_52; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_53; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_54; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_55; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_56; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_57; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_58; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_59; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_60; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_61; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_62; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_leftNodeIsCharacter_63; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_0; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_1; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_2; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_3; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_4; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_5; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_6; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_7; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_8; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_9; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_10; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_11; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_12; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_13; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_14; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_15; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_16; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_17; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_18; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_19; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_20; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_21; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_22; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_23; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_24; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_25; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_26; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_27; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_28; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_29; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_30; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_31; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_32; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_33; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_34; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_35; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_36; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_37; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_38; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_39; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_40; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_41; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_42; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_43; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_44; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_45; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_46; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_47; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_48; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_49; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_50; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_51; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_52; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_53; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_54; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_55; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_56; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_57; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_58; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_59; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_60; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_61; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_62; // @[topLevel.scala 56:18]
  wire  tg_io_outputs_rightNodeIsCharacter_63; // @[topLevel.scala 56:18]
  wire [6:0] tg_io_outputs_validNodes; // @[topLevel.scala 56:18]
  wire [5:0] tg_io_outputs_validCharacters; // @[topLevel.scala 56:18]
  wire  tg_io_finished; // @[topLevel.scala 56:18]
  wire  tdc_clock; // @[topLevel.scala 57:19]
  wire  tdc_reset; // @[topLevel.scala 57:19]
  wire  tdc_io_start; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_0; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_1; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_2; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_3; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_4; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_5; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_6; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_7; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_8; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_9; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_10; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_11; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_12; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_13; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_14; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_15; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_16; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_17; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_18; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_19; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_20; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_21; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_22; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_23; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_24; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_25; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_26; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_27; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_28; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_29; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_30; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_31; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_32; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_33; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_34; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_35; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_36; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_37; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_38; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_39; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_40; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_41; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_42; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_43; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_44; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_45; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_46; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_47; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_48; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_49; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_50; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_51; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_52; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_53; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_54; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_55; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_56; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_57; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_58; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_59; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_60; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_61; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_62; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_leftNode_63; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_0; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_1; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_2; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_3; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_4; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_5; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_6; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_7; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_8; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_9; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_10; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_11; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_12; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_13; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_14; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_15; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_16; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_17; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_18; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_19; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_20; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_21; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_22; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_23; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_24; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_25; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_26; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_27; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_28; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_29; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_30; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_31; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_32; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_33; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_34; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_35; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_36; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_37; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_38; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_39; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_40; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_41; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_42; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_43; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_44; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_45; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_46; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_47; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_48; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_49; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_50; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_51; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_52; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_53; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_54; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_55; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_56; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_57; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_58; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_59; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_60; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_61; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_62; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_inputs_rightNode_63; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_0; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_1; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_2; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_3; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_4; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_5; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_6; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_7; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_8; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_9; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_10; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_11; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_12; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_13; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_14; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_15; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_16; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_17; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_18; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_19; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_20; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_21; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_22; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_23; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_24; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_25; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_26; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_27; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_28; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_29; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_30; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_31; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_32; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_33; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_34; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_35; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_36; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_37; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_38; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_39; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_40; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_41; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_42; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_43; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_44; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_45; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_46; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_47; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_48; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_49; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_50; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_51; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_52; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_53; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_54; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_55; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_56; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_57; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_58; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_59; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_60; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_61; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_62; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_leftNodeIsCharacter_63; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_0; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_1; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_2; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_3; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_4; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_5; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_6; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_7; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_8; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_9; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_10; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_11; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_12; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_13; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_14; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_15; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_16; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_17; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_18; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_19; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_20; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_21; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_22; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_23; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_24; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_25; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_26; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_27; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_28; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_29; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_30; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_31; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_32; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_33; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_34; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_35; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_36; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_37; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_38; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_39; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_40; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_41; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_42; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_43; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_44; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_45; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_46; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_47; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_48; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_49; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_50; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_51; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_52; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_53; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_54; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_55; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_56; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_57; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_58; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_59; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_60; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_61; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_62; // @[topLevel.scala 57:19]
  wire  tdc_io_inputs_rightNodeIsCharacter_63; // @[topLevel.scala 57:19]
  wire [6:0] tdc_io_inputs_validNodes; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_inputs_validCharacters; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_0; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_1; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_2; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_3; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_4; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_5; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_6; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_7; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_8; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_9; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_10; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_11; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_12; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_13; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_14; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_15; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_16; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_17; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_18; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_19; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_20; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_21; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_22; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_23; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_24; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_25; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_26; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_27; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_28; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_29; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_30; // @[topLevel.scala 57:19]
  wire [8:0] tdc_io_outputs_characters_31; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_0; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_1; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_2; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_3; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_4; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_5; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_6; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_7; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_8; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_9; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_10; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_11; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_12; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_13; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_14; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_15; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_16; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_17; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_18; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_19; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_20; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_21; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_22; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_23; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_24; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_25; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_26; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_27; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_28; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_29; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_30; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_depths_31; // @[topLevel.scala 57:19]
  wire [5:0] tdc_io_outputs_validCharacters; // @[topLevel.scala 57:19]
  wire  tdc_io_finished; // @[topLevel.scala 57:19]
  wire  sltg_clock; // @[topLevel.scala 58:20]
  wire  sltg_reset; // @[topLevel.scala 58:20]
  wire  sltg_io_start; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_0; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_1; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_2; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_3; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_4; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_5; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_6; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_7; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_8; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_9; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_10; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_11; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_12; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_13; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_14; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_15; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_16; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_17; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_18; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_19; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_20; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_21; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_22; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_23; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_24; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_25; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_26; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_27; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_28; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_29; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_30; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_inputs_characters_31; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_0; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_1; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_2; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_3; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_4; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_5; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_6; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_7; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_8; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_9; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_10; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_11; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_12; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_13; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_14; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_15; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_16; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_17; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_18; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_19; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_20; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_21; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_22; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_23; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_24; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_25; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_26; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_27; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_28; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_29; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_30; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_depths_31; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_inputs_validCharacters; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_0; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_1; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_2; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_3; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_4; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_5; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_6; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_7; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_8; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_9; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_10; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_11; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_12; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_13; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_14; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_15; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_16; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_17; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_18; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_19; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_20; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_21; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_22; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_23; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_24; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_25; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_26; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_27; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_28; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_29; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_30; // @[topLevel.scala 58:20]
  wire [7:0] sltg_io_outputs_outputData_31; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_0; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_1; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_2; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_3; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_4; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_5; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_6; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_7; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_8; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_9; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_10; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_11; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_12; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_13; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_14; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_15; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_16; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_17; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_18; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_19; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_20; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_21; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_22; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_23; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_24; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_25; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_26; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_27; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_28; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_29; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_30; // @[topLevel.scala 58:20]
  wire [8:0] sltg_io_outputs_outputTags_31; // @[topLevel.scala 58:20]
  wire [5:0] sltg_io_outputs_itemNumber; // @[topLevel.scala 58:20]
  wire  sltg_io_finished; // @[topLevel.scala 58:20]
  wire  tn_clock; // @[topLevel.scala 59:18]
  wire  tn_reset; // @[topLevel.scala 59:18]
  wire  tn_io_start; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_0; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_1; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_2; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_3; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_4; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_5; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_6; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_7; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_8; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_9; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_10; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_11; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_12; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_13; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_14; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_15; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_16; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_17; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_18; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_19; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_20; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_21; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_22; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_23; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_24; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_25; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_26; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_27; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_28; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_29; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_30; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_inputs_outputData_31; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_0; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_1; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_2; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_3; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_4; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_5; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_6; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_7; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_8; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_9; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_10; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_11; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_12; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_13; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_14; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_15; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_16; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_17; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_18; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_19; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_20; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_21; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_22; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_23; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_24; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_25; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_26; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_27; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_28; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_29; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_30; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_inputs_outputTags_31; // @[topLevel.scala 59:18]
  wire [5:0] tn_io_inputs_itemNumber; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_0; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_1; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_2; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_3; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_4; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_5; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_6; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_7; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_8; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_9; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_10; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_11; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_12; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_13; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_14; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_15; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_16; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_17; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_18; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_19; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_20; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_21; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_22; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_23; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_24; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_25; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_26; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_27; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_28; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_29; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_30; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_charactersOut_31; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_0; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_1; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_2; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_3; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_4; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_5; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_6; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_7; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_8; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_9; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_10; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_11; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_12; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_13; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_14; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_15; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_16; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_17; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_18; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_19; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_20; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_21; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_22; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_23; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_24; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_25; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_26; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_27; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_28; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_29; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_30; // @[topLevel.scala 59:18]
  wire [7:0] tn_io_outputs_depthsOut_31; // @[topLevel.scala 59:18]
  wire [8:0] tn_io_outputs_validNodesOut; // @[topLevel.scala 59:18]
  wire  tn_io_finished; // @[topLevel.scala 59:18]
  wire  cg_clock; // @[topLevel.scala 69:18]
  wire  cg_reset; // @[topLevel.scala 69:18]
  wire  cg_io_start; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_0; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_1; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_2; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_3; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_4; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_5; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_6; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_7; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_8; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_9; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_10; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_11; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_12; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_13; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_14; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_15; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_16; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_17; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_18; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_19; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_20; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_21; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_22; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_23; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_24; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_25; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_26; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_27; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_28; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_29; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_30; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_charactersOut_31; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_0; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_1; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_2; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_3; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_4; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_5; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_6; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_7; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_8; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_9; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_10; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_11; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_12; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_13; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_14; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_15; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_16; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_17; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_18; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_19; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_20; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_21; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_22; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_23; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_24; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_25; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_26; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_27; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_28; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_29; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_30; // @[topLevel.scala 69:18]
  wire [7:0] cg_io_inputs_depthsOut_31; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_inputs_validNodesOut; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_0; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_1; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_2; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_3; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_4; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_5; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_6; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_7; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_8; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_9; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_10; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_11; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_12; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_13; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_14; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_15; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_16; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_17; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_18; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_19; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_20; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_21; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_22; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_23; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_24; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_25; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_26; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_27; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_28; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_29; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_30; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_31; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_32; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_33; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_34; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_35; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_36; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_37; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_38; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_39; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_40; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_41; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_42; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_43; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_44; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_45; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_46; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_47; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_48; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_49; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_50; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_51; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_52; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_53; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_54; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_55; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_56; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_57; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_58; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_59; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_60; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_61; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_62; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_63; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_64; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_65; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_66; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_67; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_68; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_69; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_70; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_71; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_72; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_73; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_74; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_75; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_76; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_77; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_78; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_79; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_80; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_81; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_82; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_83; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_84; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_85; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_86; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_87; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_88; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_89; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_90; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_91; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_92; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_93; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_94; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_95; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_96; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_97; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_98; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_99; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_100; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_101; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_102; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_103; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_104; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_105; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_106; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_107; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_108; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_109; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_110; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_111; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_112; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_113; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_114; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_115; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_116; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_117; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_118; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_119; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_120; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_121; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_122; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_123; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_124; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_125; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_126; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_127; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_128; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_129; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_130; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_131; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_132; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_133; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_134; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_135; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_136; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_137; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_138; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_139; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_140; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_141; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_142; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_143; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_144; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_145; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_146; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_147; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_148; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_149; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_150; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_151; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_152; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_153; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_154; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_155; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_156; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_157; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_158; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_159; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_160; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_161; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_162; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_163; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_164; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_165; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_166; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_167; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_168; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_169; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_170; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_171; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_172; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_173; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_174; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_175; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_176; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_177; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_178; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_179; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_180; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_181; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_182; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_183; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_184; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_185; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_186; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_187; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_188; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_189; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_190; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_191; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_192; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_193; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_194; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_195; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_196; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_197; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_198; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_199; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_200; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_201; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_202; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_203; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_204; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_205; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_206; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_207; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_208; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_209; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_210; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_211; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_212; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_213; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_214; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_215; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_216; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_217; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_218; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_219; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_220; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_221; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_222; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_223; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_224; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_225; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_226; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_227; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_228; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_229; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_230; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_231; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_232; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_233; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_234; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_235; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_236; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_237; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_238; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_239; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_240; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_241; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_242; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_243; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_244; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_245; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_246; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_247; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_248; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_249; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_250; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_251; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_252; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_253; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_254; // @[topLevel.scala 69:18]
  wire [23:0] cg_io_outputs_codewords_255; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_0; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_1; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_2; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_3; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_4; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_5; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_6; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_7; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_8; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_9; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_10; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_11; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_12; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_13; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_14; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_15; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_16; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_17; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_18; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_19; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_20; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_21; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_22; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_23; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_24; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_25; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_26; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_27; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_28; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_29; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_30; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_31; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_32; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_33; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_34; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_35; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_36; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_37; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_38; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_39; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_40; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_41; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_42; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_43; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_44; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_45; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_46; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_47; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_48; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_49; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_50; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_51; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_52; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_53; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_54; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_55; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_56; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_57; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_58; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_59; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_60; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_61; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_62; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_63; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_64; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_65; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_66; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_67; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_68; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_69; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_70; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_71; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_72; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_73; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_74; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_75; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_76; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_77; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_78; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_79; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_80; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_81; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_82; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_83; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_84; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_85; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_86; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_87; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_88; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_89; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_90; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_91; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_92; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_93; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_94; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_95; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_96; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_97; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_98; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_99; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_100; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_101; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_102; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_103; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_104; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_105; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_106; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_107; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_108; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_109; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_110; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_111; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_112; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_113; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_114; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_115; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_116; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_117; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_118; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_119; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_120; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_121; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_122; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_123; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_124; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_125; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_126; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_127; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_128; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_129; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_130; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_131; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_132; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_133; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_134; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_135; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_136; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_137; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_138; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_139; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_140; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_141; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_142; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_143; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_144; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_145; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_146; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_147; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_148; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_149; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_150; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_151; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_152; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_153; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_154; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_155; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_156; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_157; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_158; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_159; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_160; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_161; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_162; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_163; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_164; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_165; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_166; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_167; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_168; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_169; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_170; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_171; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_172; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_173; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_174; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_175; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_176; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_177; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_178; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_179; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_180; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_181; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_182; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_183; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_184; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_185; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_186; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_187; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_188; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_189; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_190; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_191; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_192; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_193; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_194; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_195; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_196; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_197; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_198; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_199; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_200; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_201; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_202; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_203; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_204; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_205; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_206; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_207; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_208; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_209; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_210; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_211; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_212; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_213; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_214; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_215; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_216; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_217; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_218; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_219; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_220; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_221; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_222; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_223; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_224; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_225; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_226; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_227; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_228; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_229; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_230; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_231; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_232; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_233; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_234; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_235; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_236; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_237; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_238; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_239; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_240; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_241; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_242; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_243; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_244; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_245; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_246; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_247; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_248; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_249; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_250; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_251; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_252; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_253; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_254; // @[topLevel.scala 69:18]
  wire [4:0] cg_io_outputs_lengths_255; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_0; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_1; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_2; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_3; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_4; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_5; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_6; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_7; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_8; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_9; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_10; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_11; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_12; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_13; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_14; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_15; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_16; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_17; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_18; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_19; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_20; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_21; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_22; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_23; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_24; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_25; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_26; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_27; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_28; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_29; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_30; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_charactersOut_31; // @[topLevel.scala 69:18]
  wire [8:0] cg_io_outputs_nodes; // @[topLevel.scala 69:18]
  wire [3:0] cg_io_outputs_escapeCharacterLength; // @[topLevel.scala 69:18]
  wire [15:0] cg_io_outputs_escapeCodeword; // @[topLevel.scala 69:18]
  wire  cg_io_finished; // @[topLevel.scala 69:18]
  wire  co_clock; // @[topLevel.scala 72:18]
  wire  co_reset; // @[topLevel.scala 72:18]
  wire  co_io_start; // @[topLevel.scala 72:18]
  wire [11:0] co_io_dataIn_0_currentByteOut; // @[topLevel.scala 72:18]
  wire [7:0] co_io_dataIn_0_dataIn_0; // @[topLevel.scala 72:18]
  wire  co_io_dataIn_0_valid; // @[topLevel.scala 72:18]
  wire  co_io_dataIn_0_ready; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_0; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_1; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_2; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_3; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_4; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_5; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_6; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_7; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_8; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_9; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_10; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_11; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_12; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_13; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_14; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_15; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_16; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_17; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_18; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_19; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_20; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_21; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_22; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_23; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_24; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_25; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_26; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_27; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_28; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_29; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_30; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_31; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_32; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_33; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_34; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_35; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_36; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_37; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_38; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_39; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_40; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_41; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_42; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_43; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_44; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_45; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_46; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_47; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_48; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_49; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_50; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_51; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_52; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_53; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_54; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_55; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_56; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_57; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_58; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_59; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_60; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_61; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_62; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_63; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_64; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_65; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_66; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_67; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_68; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_69; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_70; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_71; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_72; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_73; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_74; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_75; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_76; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_77; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_78; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_79; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_80; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_81; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_82; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_83; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_84; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_85; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_86; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_87; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_88; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_89; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_90; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_91; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_92; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_93; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_94; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_95; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_96; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_97; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_98; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_99; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_100; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_101; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_102; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_103; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_104; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_105; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_106; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_107; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_108; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_109; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_110; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_111; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_112; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_113; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_114; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_115; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_116; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_117; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_118; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_119; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_120; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_121; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_122; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_123; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_124; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_125; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_126; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_127; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_128; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_129; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_130; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_131; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_132; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_133; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_134; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_135; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_136; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_137; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_138; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_139; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_140; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_141; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_142; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_143; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_144; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_145; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_146; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_147; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_148; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_149; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_150; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_151; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_152; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_153; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_154; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_155; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_156; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_157; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_158; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_159; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_160; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_161; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_162; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_163; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_164; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_165; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_166; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_167; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_168; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_169; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_170; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_171; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_172; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_173; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_174; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_175; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_176; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_177; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_178; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_179; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_180; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_181; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_182; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_183; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_184; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_185; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_186; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_187; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_188; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_189; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_190; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_191; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_192; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_193; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_194; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_195; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_196; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_197; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_198; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_199; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_200; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_201; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_202; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_203; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_204; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_205; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_206; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_207; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_208; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_209; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_210; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_211; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_212; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_213; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_214; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_215; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_216; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_217; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_218; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_219; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_220; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_221; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_222; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_223; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_224; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_225; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_226; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_227; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_228; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_229; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_230; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_231; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_232; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_233; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_234; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_235; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_236; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_237; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_238; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_239; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_240; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_241; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_242; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_243; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_244; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_245; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_246; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_247; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_248; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_249; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_250; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_251; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_252; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_253; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_254; // @[topLevel.scala 72:18]
  wire [23:0] co_io_inputs_codewords_255; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_0; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_1; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_2; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_3; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_4; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_5; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_6; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_7; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_8; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_9; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_10; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_11; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_12; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_13; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_14; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_15; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_16; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_17; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_18; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_19; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_20; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_21; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_22; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_23; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_24; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_25; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_26; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_27; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_28; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_29; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_30; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_31; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_32; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_33; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_34; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_35; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_36; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_37; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_38; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_39; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_40; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_41; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_42; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_43; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_44; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_45; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_46; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_47; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_48; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_49; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_50; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_51; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_52; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_53; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_54; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_55; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_56; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_57; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_58; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_59; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_60; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_61; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_62; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_63; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_64; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_65; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_66; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_67; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_68; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_69; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_70; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_71; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_72; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_73; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_74; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_75; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_76; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_77; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_78; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_79; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_80; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_81; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_82; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_83; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_84; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_85; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_86; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_87; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_88; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_89; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_90; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_91; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_92; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_93; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_94; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_95; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_96; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_97; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_98; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_99; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_100; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_101; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_102; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_103; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_104; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_105; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_106; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_107; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_108; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_109; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_110; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_111; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_112; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_113; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_114; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_115; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_116; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_117; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_118; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_119; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_120; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_121; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_122; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_123; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_124; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_125; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_126; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_127; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_128; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_129; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_130; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_131; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_132; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_133; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_134; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_135; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_136; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_137; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_138; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_139; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_140; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_141; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_142; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_143; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_144; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_145; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_146; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_147; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_148; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_149; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_150; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_151; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_152; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_153; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_154; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_155; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_156; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_157; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_158; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_159; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_160; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_161; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_162; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_163; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_164; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_165; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_166; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_167; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_168; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_169; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_170; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_171; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_172; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_173; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_174; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_175; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_176; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_177; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_178; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_179; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_180; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_181; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_182; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_183; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_184; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_185; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_186; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_187; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_188; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_189; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_190; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_191; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_192; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_193; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_194; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_195; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_196; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_197; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_198; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_199; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_200; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_201; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_202; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_203; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_204; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_205; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_206; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_207; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_208; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_209; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_210; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_211; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_212; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_213; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_214; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_215; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_216; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_217; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_218; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_219; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_220; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_221; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_222; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_223; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_224; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_225; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_226; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_227; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_228; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_229; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_230; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_231; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_232; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_233; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_234; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_235; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_236; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_237; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_238; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_239; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_240; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_241; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_242; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_243; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_244; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_245; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_246; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_247; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_248; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_249; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_250; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_251; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_252; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_253; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_254; // @[topLevel.scala 72:18]
  wire [4:0] co_io_inputs_lengths_255; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_0; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_1; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_2; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_3; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_4; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_5; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_6; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_7; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_8; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_9; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_10; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_11; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_12; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_13; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_14; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_15; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_16; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_17; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_18; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_19; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_20; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_21; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_22; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_23; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_24; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_25; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_26; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_27; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_28; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_29; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_30; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_charactersOut_31; // @[topLevel.scala 72:18]
  wire [8:0] co_io_inputs_nodes; // @[topLevel.scala 72:18]
  wire [3:0] co_io_inputs_escapeCharacterLength; // @[topLevel.scala 72:18]
  wire [15:0] co_io_inputs_escapeCodeword; // @[topLevel.scala 72:18]
  wire [27:0] co_io_outputs_0_dataOut; // @[topLevel.scala 72:18]
  wire [4:0] co_io_outputs_0_dataLength; // @[topLevel.scala 72:18]
  wire  co_io_outputs_0_valid; // @[topLevel.scala 72:18]
  wire  co_io_outputs_0_ready; // @[topLevel.scala 72:18]
  wire  co_io_finished; // @[topLevel.scala 72:18]
  reg  previousStart; // @[topLevel.scala 75:30]
  reg [31:0] _RAND_0;
  reg  cfmPreviousFinished; // @[topLevel.scala 76:36]
  reg [31:0] _RAND_1;
  reg  tgPreviousFinished; // @[topLevel.scala 77:35]
  reg [31:0] _RAND_2;
  reg  tdcPreviousFinished; // @[topLevel.scala 78:36]
  reg [31:0] _RAND_3;
  reg  sltgPreviousFinished; // @[topLevel.scala 79:37]
  reg [31:0] _RAND_4;
  reg  tnPreviousFinished; // @[topLevel.scala 80:35]
  reg [31:0] _RAND_5;
  reg  cgPreviousFinished; // @[topLevel.scala 81:35]
  reg [31:0] _RAND_6;
  reg  coPreviousFinished; // @[topLevel.scala 82:35]
  reg [31:0] _RAND_7;
  wire  _T = ~previousStart; // @[topLevel.scala 83:31]
  wire  _T_2 = ~cfmPreviousFinished; // @[topLevel.scala 84:37]
  wire  _T_4 = ~tgPreviousFinished; // @[topLevel.scala 85:37]
  wire  _T_6 = ~tdcPreviousFinished; // @[topLevel.scala 86:39]
  wire  _T_8 = ~sltgPreviousFinished; // @[topLevel.scala 87:38]
  wire  _T_10 = ~tnPreviousFinished; // @[topLevel.scala 88:36]
  wire  _T_12 = ~cgPreviousFinished; // @[topLevel.scala 89:36]
  wire  _T_14 = ~coPreviousFinished; // @[topLevel.scala 90:36]
  characterFrequencyModule cfm ( // @[topLevel.scala 55:19]
    .clock(cfm_clock),
    .reset(cfm_reset),
    .io_start(cfm_io_start),
    .io_input_currentByteOut(cfm_io_input_currentByteOut),
    .io_input_dataIn_0(cfm_io_input_dataIn_0),
    .io_input_valid(cfm_io_input_valid),
    .io_input_ready(cfm_io_input_ready),
    .io_outputs_sortedFrequency_0(cfm_io_outputs_sortedFrequency_0),
    .io_outputs_sortedFrequency_1(cfm_io_outputs_sortedFrequency_1),
    .io_outputs_sortedFrequency_2(cfm_io_outputs_sortedFrequency_2),
    .io_outputs_sortedFrequency_3(cfm_io_outputs_sortedFrequency_3),
    .io_outputs_sortedFrequency_4(cfm_io_outputs_sortedFrequency_4),
    .io_outputs_sortedFrequency_5(cfm_io_outputs_sortedFrequency_5),
    .io_outputs_sortedFrequency_6(cfm_io_outputs_sortedFrequency_6),
    .io_outputs_sortedFrequency_7(cfm_io_outputs_sortedFrequency_7),
    .io_outputs_sortedFrequency_8(cfm_io_outputs_sortedFrequency_8),
    .io_outputs_sortedFrequency_9(cfm_io_outputs_sortedFrequency_9),
    .io_outputs_sortedFrequency_10(cfm_io_outputs_sortedFrequency_10),
    .io_outputs_sortedFrequency_11(cfm_io_outputs_sortedFrequency_11),
    .io_outputs_sortedFrequency_12(cfm_io_outputs_sortedFrequency_12),
    .io_outputs_sortedFrequency_13(cfm_io_outputs_sortedFrequency_13),
    .io_outputs_sortedFrequency_14(cfm_io_outputs_sortedFrequency_14),
    .io_outputs_sortedFrequency_15(cfm_io_outputs_sortedFrequency_15),
    .io_outputs_sortedFrequency_16(cfm_io_outputs_sortedFrequency_16),
    .io_outputs_sortedFrequency_17(cfm_io_outputs_sortedFrequency_17),
    .io_outputs_sortedFrequency_18(cfm_io_outputs_sortedFrequency_18),
    .io_outputs_sortedFrequency_19(cfm_io_outputs_sortedFrequency_19),
    .io_outputs_sortedFrequency_20(cfm_io_outputs_sortedFrequency_20),
    .io_outputs_sortedFrequency_21(cfm_io_outputs_sortedFrequency_21),
    .io_outputs_sortedFrequency_22(cfm_io_outputs_sortedFrequency_22),
    .io_outputs_sortedFrequency_23(cfm_io_outputs_sortedFrequency_23),
    .io_outputs_sortedFrequency_24(cfm_io_outputs_sortedFrequency_24),
    .io_outputs_sortedFrequency_25(cfm_io_outputs_sortedFrequency_25),
    .io_outputs_sortedFrequency_26(cfm_io_outputs_sortedFrequency_26),
    .io_outputs_sortedFrequency_27(cfm_io_outputs_sortedFrequency_27),
    .io_outputs_sortedFrequency_28(cfm_io_outputs_sortedFrequency_28),
    .io_outputs_sortedFrequency_29(cfm_io_outputs_sortedFrequency_29),
    .io_outputs_sortedFrequency_30(cfm_io_outputs_sortedFrequency_30),
    .io_outputs_sortedFrequency_31(cfm_io_outputs_sortedFrequency_31),
    .io_outputs_sortedCharacter_0(cfm_io_outputs_sortedCharacter_0),
    .io_outputs_sortedCharacter_1(cfm_io_outputs_sortedCharacter_1),
    .io_outputs_sortedCharacter_2(cfm_io_outputs_sortedCharacter_2),
    .io_outputs_sortedCharacter_3(cfm_io_outputs_sortedCharacter_3),
    .io_outputs_sortedCharacter_4(cfm_io_outputs_sortedCharacter_4),
    .io_outputs_sortedCharacter_5(cfm_io_outputs_sortedCharacter_5),
    .io_outputs_sortedCharacter_6(cfm_io_outputs_sortedCharacter_6),
    .io_outputs_sortedCharacter_7(cfm_io_outputs_sortedCharacter_7),
    .io_outputs_sortedCharacter_8(cfm_io_outputs_sortedCharacter_8),
    .io_outputs_sortedCharacter_9(cfm_io_outputs_sortedCharacter_9),
    .io_outputs_sortedCharacter_10(cfm_io_outputs_sortedCharacter_10),
    .io_outputs_sortedCharacter_11(cfm_io_outputs_sortedCharacter_11),
    .io_outputs_sortedCharacter_12(cfm_io_outputs_sortedCharacter_12),
    .io_outputs_sortedCharacter_13(cfm_io_outputs_sortedCharacter_13),
    .io_outputs_sortedCharacter_14(cfm_io_outputs_sortedCharacter_14),
    .io_outputs_sortedCharacter_15(cfm_io_outputs_sortedCharacter_15),
    .io_outputs_sortedCharacter_16(cfm_io_outputs_sortedCharacter_16),
    .io_outputs_sortedCharacter_17(cfm_io_outputs_sortedCharacter_17),
    .io_outputs_sortedCharacter_18(cfm_io_outputs_sortedCharacter_18),
    .io_outputs_sortedCharacter_19(cfm_io_outputs_sortedCharacter_19),
    .io_outputs_sortedCharacter_20(cfm_io_outputs_sortedCharacter_20),
    .io_outputs_sortedCharacter_21(cfm_io_outputs_sortedCharacter_21),
    .io_outputs_sortedCharacter_22(cfm_io_outputs_sortedCharacter_22),
    .io_outputs_sortedCharacter_23(cfm_io_outputs_sortedCharacter_23),
    .io_outputs_sortedCharacter_24(cfm_io_outputs_sortedCharacter_24),
    .io_outputs_sortedCharacter_25(cfm_io_outputs_sortedCharacter_25),
    .io_outputs_sortedCharacter_26(cfm_io_outputs_sortedCharacter_26),
    .io_outputs_sortedCharacter_27(cfm_io_outputs_sortedCharacter_27),
    .io_outputs_sortedCharacter_28(cfm_io_outputs_sortedCharacter_28),
    .io_outputs_sortedCharacter_29(cfm_io_outputs_sortedCharacter_29),
    .io_outputs_sortedCharacter_30(cfm_io_outputs_sortedCharacter_30),
    .io_outputs_sortedCharacter_31(cfm_io_outputs_sortedCharacter_31),
    .io_finished(cfm_io_finished)
  );
  treeGenerator tg ( // @[topLevel.scala 56:18]
    .clock(tg_clock),
    .reset(tg_reset),
    .io_start(tg_io_start),
    .io_inputs_sortedFrequency_0(tg_io_inputs_sortedFrequency_0),
    .io_inputs_sortedFrequency_1(tg_io_inputs_sortedFrequency_1),
    .io_inputs_sortedFrequency_2(tg_io_inputs_sortedFrequency_2),
    .io_inputs_sortedFrequency_3(tg_io_inputs_sortedFrequency_3),
    .io_inputs_sortedFrequency_4(tg_io_inputs_sortedFrequency_4),
    .io_inputs_sortedFrequency_5(tg_io_inputs_sortedFrequency_5),
    .io_inputs_sortedFrequency_6(tg_io_inputs_sortedFrequency_6),
    .io_inputs_sortedFrequency_7(tg_io_inputs_sortedFrequency_7),
    .io_inputs_sortedFrequency_8(tg_io_inputs_sortedFrequency_8),
    .io_inputs_sortedFrequency_9(tg_io_inputs_sortedFrequency_9),
    .io_inputs_sortedFrequency_10(tg_io_inputs_sortedFrequency_10),
    .io_inputs_sortedFrequency_11(tg_io_inputs_sortedFrequency_11),
    .io_inputs_sortedFrequency_12(tg_io_inputs_sortedFrequency_12),
    .io_inputs_sortedFrequency_13(tg_io_inputs_sortedFrequency_13),
    .io_inputs_sortedFrequency_14(tg_io_inputs_sortedFrequency_14),
    .io_inputs_sortedFrequency_15(tg_io_inputs_sortedFrequency_15),
    .io_inputs_sortedFrequency_16(tg_io_inputs_sortedFrequency_16),
    .io_inputs_sortedFrequency_17(tg_io_inputs_sortedFrequency_17),
    .io_inputs_sortedFrequency_18(tg_io_inputs_sortedFrequency_18),
    .io_inputs_sortedFrequency_19(tg_io_inputs_sortedFrequency_19),
    .io_inputs_sortedFrequency_20(tg_io_inputs_sortedFrequency_20),
    .io_inputs_sortedFrequency_21(tg_io_inputs_sortedFrequency_21),
    .io_inputs_sortedFrequency_22(tg_io_inputs_sortedFrequency_22),
    .io_inputs_sortedFrequency_23(tg_io_inputs_sortedFrequency_23),
    .io_inputs_sortedFrequency_24(tg_io_inputs_sortedFrequency_24),
    .io_inputs_sortedFrequency_25(tg_io_inputs_sortedFrequency_25),
    .io_inputs_sortedFrequency_26(tg_io_inputs_sortedFrequency_26),
    .io_inputs_sortedFrequency_27(tg_io_inputs_sortedFrequency_27),
    .io_inputs_sortedFrequency_28(tg_io_inputs_sortedFrequency_28),
    .io_inputs_sortedFrequency_29(tg_io_inputs_sortedFrequency_29),
    .io_inputs_sortedFrequency_30(tg_io_inputs_sortedFrequency_30),
    .io_inputs_sortedFrequency_31(tg_io_inputs_sortedFrequency_31),
    .io_inputs_sortedCharacter_0(tg_io_inputs_sortedCharacter_0),
    .io_inputs_sortedCharacter_1(tg_io_inputs_sortedCharacter_1),
    .io_inputs_sortedCharacter_2(tg_io_inputs_sortedCharacter_2),
    .io_inputs_sortedCharacter_3(tg_io_inputs_sortedCharacter_3),
    .io_inputs_sortedCharacter_4(tg_io_inputs_sortedCharacter_4),
    .io_inputs_sortedCharacter_5(tg_io_inputs_sortedCharacter_5),
    .io_inputs_sortedCharacter_6(tg_io_inputs_sortedCharacter_6),
    .io_inputs_sortedCharacter_7(tg_io_inputs_sortedCharacter_7),
    .io_inputs_sortedCharacter_8(tg_io_inputs_sortedCharacter_8),
    .io_inputs_sortedCharacter_9(tg_io_inputs_sortedCharacter_9),
    .io_inputs_sortedCharacter_10(tg_io_inputs_sortedCharacter_10),
    .io_inputs_sortedCharacter_11(tg_io_inputs_sortedCharacter_11),
    .io_inputs_sortedCharacter_12(tg_io_inputs_sortedCharacter_12),
    .io_inputs_sortedCharacter_13(tg_io_inputs_sortedCharacter_13),
    .io_inputs_sortedCharacter_14(tg_io_inputs_sortedCharacter_14),
    .io_inputs_sortedCharacter_15(tg_io_inputs_sortedCharacter_15),
    .io_inputs_sortedCharacter_16(tg_io_inputs_sortedCharacter_16),
    .io_inputs_sortedCharacter_17(tg_io_inputs_sortedCharacter_17),
    .io_inputs_sortedCharacter_18(tg_io_inputs_sortedCharacter_18),
    .io_inputs_sortedCharacter_19(tg_io_inputs_sortedCharacter_19),
    .io_inputs_sortedCharacter_20(tg_io_inputs_sortedCharacter_20),
    .io_inputs_sortedCharacter_21(tg_io_inputs_sortedCharacter_21),
    .io_inputs_sortedCharacter_22(tg_io_inputs_sortedCharacter_22),
    .io_inputs_sortedCharacter_23(tg_io_inputs_sortedCharacter_23),
    .io_inputs_sortedCharacter_24(tg_io_inputs_sortedCharacter_24),
    .io_inputs_sortedCharacter_25(tg_io_inputs_sortedCharacter_25),
    .io_inputs_sortedCharacter_26(tg_io_inputs_sortedCharacter_26),
    .io_inputs_sortedCharacter_27(tg_io_inputs_sortedCharacter_27),
    .io_inputs_sortedCharacter_28(tg_io_inputs_sortedCharacter_28),
    .io_inputs_sortedCharacter_29(tg_io_inputs_sortedCharacter_29),
    .io_inputs_sortedCharacter_30(tg_io_inputs_sortedCharacter_30),
    .io_inputs_sortedCharacter_31(tg_io_inputs_sortedCharacter_31),
    .io_outputs_leftNode_0(tg_io_outputs_leftNode_0),
    .io_outputs_leftNode_1(tg_io_outputs_leftNode_1),
    .io_outputs_leftNode_2(tg_io_outputs_leftNode_2),
    .io_outputs_leftNode_3(tg_io_outputs_leftNode_3),
    .io_outputs_leftNode_4(tg_io_outputs_leftNode_4),
    .io_outputs_leftNode_5(tg_io_outputs_leftNode_5),
    .io_outputs_leftNode_6(tg_io_outputs_leftNode_6),
    .io_outputs_leftNode_7(tg_io_outputs_leftNode_7),
    .io_outputs_leftNode_8(tg_io_outputs_leftNode_8),
    .io_outputs_leftNode_9(tg_io_outputs_leftNode_9),
    .io_outputs_leftNode_10(tg_io_outputs_leftNode_10),
    .io_outputs_leftNode_11(tg_io_outputs_leftNode_11),
    .io_outputs_leftNode_12(tg_io_outputs_leftNode_12),
    .io_outputs_leftNode_13(tg_io_outputs_leftNode_13),
    .io_outputs_leftNode_14(tg_io_outputs_leftNode_14),
    .io_outputs_leftNode_15(tg_io_outputs_leftNode_15),
    .io_outputs_leftNode_16(tg_io_outputs_leftNode_16),
    .io_outputs_leftNode_17(tg_io_outputs_leftNode_17),
    .io_outputs_leftNode_18(tg_io_outputs_leftNode_18),
    .io_outputs_leftNode_19(tg_io_outputs_leftNode_19),
    .io_outputs_leftNode_20(tg_io_outputs_leftNode_20),
    .io_outputs_leftNode_21(tg_io_outputs_leftNode_21),
    .io_outputs_leftNode_22(tg_io_outputs_leftNode_22),
    .io_outputs_leftNode_23(tg_io_outputs_leftNode_23),
    .io_outputs_leftNode_24(tg_io_outputs_leftNode_24),
    .io_outputs_leftNode_25(tg_io_outputs_leftNode_25),
    .io_outputs_leftNode_26(tg_io_outputs_leftNode_26),
    .io_outputs_leftNode_27(tg_io_outputs_leftNode_27),
    .io_outputs_leftNode_28(tg_io_outputs_leftNode_28),
    .io_outputs_leftNode_29(tg_io_outputs_leftNode_29),
    .io_outputs_leftNode_30(tg_io_outputs_leftNode_30),
    .io_outputs_leftNode_31(tg_io_outputs_leftNode_31),
    .io_outputs_leftNode_32(tg_io_outputs_leftNode_32),
    .io_outputs_leftNode_33(tg_io_outputs_leftNode_33),
    .io_outputs_leftNode_34(tg_io_outputs_leftNode_34),
    .io_outputs_leftNode_35(tg_io_outputs_leftNode_35),
    .io_outputs_leftNode_36(tg_io_outputs_leftNode_36),
    .io_outputs_leftNode_37(tg_io_outputs_leftNode_37),
    .io_outputs_leftNode_38(tg_io_outputs_leftNode_38),
    .io_outputs_leftNode_39(tg_io_outputs_leftNode_39),
    .io_outputs_leftNode_40(tg_io_outputs_leftNode_40),
    .io_outputs_leftNode_41(tg_io_outputs_leftNode_41),
    .io_outputs_leftNode_42(tg_io_outputs_leftNode_42),
    .io_outputs_leftNode_43(tg_io_outputs_leftNode_43),
    .io_outputs_leftNode_44(tg_io_outputs_leftNode_44),
    .io_outputs_leftNode_45(tg_io_outputs_leftNode_45),
    .io_outputs_leftNode_46(tg_io_outputs_leftNode_46),
    .io_outputs_leftNode_47(tg_io_outputs_leftNode_47),
    .io_outputs_leftNode_48(tg_io_outputs_leftNode_48),
    .io_outputs_leftNode_49(tg_io_outputs_leftNode_49),
    .io_outputs_leftNode_50(tg_io_outputs_leftNode_50),
    .io_outputs_leftNode_51(tg_io_outputs_leftNode_51),
    .io_outputs_leftNode_52(tg_io_outputs_leftNode_52),
    .io_outputs_leftNode_53(tg_io_outputs_leftNode_53),
    .io_outputs_leftNode_54(tg_io_outputs_leftNode_54),
    .io_outputs_leftNode_55(tg_io_outputs_leftNode_55),
    .io_outputs_leftNode_56(tg_io_outputs_leftNode_56),
    .io_outputs_leftNode_57(tg_io_outputs_leftNode_57),
    .io_outputs_leftNode_58(tg_io_outputs_leftNode_58),
    .io_outputs_leftNode_59(tg_io_outputs_leftNode_59),
    .io_outputs_leftNode_60(tg_io_outputs_leftNode_60),
    .io_outputs_leftNode_61(tg_io_outputs_leftNode_61),
    .io_outputs_leftNode_62(tg_io_outputs_leftNode_62),
    .io_outputs_leftNode_63(tg_io_outputs_leftNode_63),
    .io_outputs_rightNode_0(tg_io_outputs_rightNode_0),
    .io_outputs_rightNode_1(tg_io_outputs_rightNode_1),
    .io_outputs_rightNode_2(tg_io_outputs_rightNode_2),
    .io_outputs_rightNode_3(tg_io_outputs_rightNode_3),
    .io_outputs_rightNode_4(tg_io_outputs_rightNode_4),
    .io_outputs_rightNode_5(tg_io_outputs_rightNode_5),
    .io_outputs_rightNode_6(tg_io_outputs_rightNode_6),
    .io_outputs_rightNode_7(tg_io_outputs_rightNode_7),
    .io_outputs_rightNode_8(tg_io_outputs_rightNode_8),
    .io_outputs_rightNode_9(tg_io_outputs_rightNode_9),
    .io_outputs_rightNode_10(tg_io_outputs_rightNode_10),
    .io_outputs_rightNode_11(tg_io_outputs_rightNode_11),
    .io_outputs_rightNode_12(tg_io_outputs_rightNode_12),
    .io_outputs_rightNode_13(tg_io_outputs_rightNode_13),
    .io_outputs_rightNode_14(tg_io_outputs_rightNode_14),
    .io_outputs_rightNode_15(tg_io_outputs_rightNode_15),
    .io_outputs_rightNode_16(tg_io_outputs_rightNode_16),
    .io_outputs_rightNode_17(tg_io_outputs_rightNode_17),
    .io_outputs_rightNode_18(tg_io_outputs_rightNode_18),
    .io_outputs_rightNode_19(tg_io_outputs_rightNode_19),
    .io_outputs_rightNode_20(tg_io_outputs_rightNode_20),
    .io_outputs_rightNode_21(tg_io_outputs_rightNode_21),
    .io_outputs_rightNode_22(tg_io_outputs_rightNode_22),
    .io_outputs_rightNode_23(tg_io_outputs_rightNode_23),
    .io_outputs_rightNode_24(tg_io_outputs_rightNode_24),
    .io_outputs_rightNode_25(tg_io_outputs_rightNode_25),
    .io_outputs_rightNode_26(tg_io_outputs_rightNode_26),
    .io_outputs_rightNode_27(tg_io_outputs_rightNode_27),
    .io_outputs_rightNode_28(tg_io_outputs_rightNode_28),
    .io_outputs_rightNode_29(tg_io_outputs_rightNode_29),
    .io_outputs_rightNode_30(tg_io_outputs_rightNode_30),
    .io_outputs_rightNode_31(tg_io_outputs_rightNode_31),
    .io_outputs_rightNode_32(tg_io_outputs_rightNode_32),
    .io_outputs_rightNode_33(tg_io_outputs_rightNode_33),
    .io_outputs_rightNode_34(tg_io_outputs_rightNode_34),
    .io_outputs_rightNode_35(tg_io_outputs_rightNode_35),
    .io_outputs_rightNode_36(tg_io_outputs_rightNode_36),
    .io_outputs_rightNode_37(tg_io_outputs_rightNode_37),
    .io_outputs_rightNode_38(tg_io_outputs_rightNode_38),
    .io_outputs_rightNode_39(tg_io_outputs_rightNode_39),
    .io_outputs_rightNode_40(tg_io_outputs_rightNode_40),
    .io_outputs_rightNode_41(tg_io_outputs_rightNode_41),
    .io_outputs_rightNode_42(tg_io_outputs_rightNode_42),
    .io_outputs_rightNode_43(tg_io_outputs_rightNode_43),
    .io_outputs_rightNode_44(tg_io_outputs_rightNode_44),
    .io_outputs_rightNode_45(tg_io_outputs_rightNode_45),
    .io_outputs_rightNode_46(tg_io_outputs_rightNode_46),
    .io_outputs_rightNode_47(tg_io_outputs_rightNode_47),
    .io_outputs_rightNode_48(tg_io_outputs_rightNode_48),
    .io_outputs_rightNode_49(tg_io_outputs_rightNode_49),
    .io_outputs_rightNode_50(tg_io_outputs_rightNode_50),
    .io_outputs_rightNode_51(tg_io_outputs_rightNode_51),
    .io_outputs_rightNode_52(tg_io_outputs_rightNode_52),
    .io_outputs_rightNode_53(tg_io_outputs_rightNode_53),
    .io_outputs_rightNode_54(tg_io_outputs_rightNode_54),
    .io_outputs_rightNode_55(tg_io_outputs_rightNode_55),
    .io_outputs_rightNode_56(tg_io_outputs_rightNode_56),
    .io_outputs_rightNode_57(tg_io_outputs_rightNode_57),
    .io_outputs_rightNode_58(tg_io_outputs_rightNode_58),
    .io_outputs_rightNode_59(tg_io_outputs_rightNode_59),
    .io_outputs_rightNode_60(tg_io_outputs_rightNode_60),
    .io_outputs_rightNode_61(tg_io_outputs_rightNode_61),
    .io_outputs_rightNode_62(tg_io_outputs_rightNode_62),
    .io_outputs_rightNode_63(tg_io_outputs_rightNode_63),
    .io_outputs_leftNodeIsCharacter_0(tg_io_outputs_leftNodeIsCharacter_0),
    .io_outputs_leftNodeIsCharacter_1(tg_io_outputs_leftNodeIsCharacter_1),
    .io_outputs_leftNodeIsCharacter_2(tg_io_outputs_leftNodeIsCharacter_2),
    .io_outputs_leftNodeIsCharacter_3(tg_io_outputs_leftNodeIsCharacter_3),
    .io_outputs_leftNodeIsCharacter_4(tg_io_outputs_leftNodeIsCharacter_4),
    .io_outputs_leftNodeIsCharacter_5(tg_io_outputs_leftNodeIsCharacter_5),
    .io_outputs_leftNodeIsCharacter_6(tg_io_outputs_leftNodeIsCharacter_6),
    .io_outputs_leftNodeIsCharacter_7(tg_io_outputs_leftNodeIsCharacter_7),
    .io_outputs_leftNodeIsCharacter_8(tg_io_outputs_leftNodeIsCharacter_8),
    .io_outputs_leftNodeIsCharacter_9(tg_io_outputs_leftNodeIsCharacter_9),
    .io_outputs_leftNodeIsCharacter_10(tg_io_outputs_leftNodeIsCharacter_10),
    .io_outputs_leftNodeIsCharacter_11(tg_io_outputs_leftNodeIsCharacter_11),
    .io_outputs_leftNodeIsCharacter_12(tg_io_outputs_leftNodeIsCharacter_12),
    .io_outputs_leftNodeIsCharacter_13(tg_io_outputs_leftNodeIsCharacter_13),
    .io_outputs_leftNodeIsCharacter_14(tg_io_outputs_leftNodeIsCharacter_14),
    .io_outputs_leftNodeIsCharacter_15(tg_io_outputs_leftNodeIsCharacter_15),
    .io_outputs_leftNodeIsCharacter_16(tg_io_outputs_leftNodeIsCharacter_16),
    .io_outputs_leftNodeIsCharacter_17(tg_io_outputs_leftNodeIsCharacter_17),
    .io_outputs_leftNodeIsCharacter_18(tg_io_outputs_leftNodeIsCharacter_18),
    .io_outputs_leftNodeIsCharacter_19(tg_io_outputs_leftNodeIsCharacter_19),
    .io_outputs_leftNodeIsCharacter_20(tg_io_outputs_leftNodeIsCharacter_20),
    .io_outputs_leftNodeIsCharacter_21(tg_io_outputs_leftNodeIsCharacter_21),
    .io_outputs_leftNodeIsCharacter_22(tg_io_outputs_leftNodeIsCharacter_22),
    .io_outputs_leftNodeIsCharacter_23(tg_io_outputs_leftNodeIsCharacter_23),
    .io_outputs_leftNodeIsCharacter_24(tg_io_outputs_leftNodeIsCharacter_24),
    .io_outputs_leftNodeIsCharacter_25(tg_io_outputs_leftNodeIsCharacter_25),
    .io_outputs_leftNodeIsCharacter_26(tg_io_outputs_leftNodeIsCharacter_26),
    .io_outputs_leftNodeIsCharacter_27(tg_io_outputs_leftNodeIsCharacter_27),
    .io_outputs_leftNodeIsCharacter_28(tg_io_outputs_leftNodeIsCharacter_28),
    .io_outputs_leftNodeIsCharacter_29(tg_io_outputs_leftNodeIsCharacter_29),
    .io_outputs_leftNodeIsCharacter_30(tg_io_outputs_leftNodeIsCharacter_30),
    .io_outputs_leftNodeIsCharacter_31(tg_io_outputs_leftNodeIsCharacter_31),
    .io_outputs_leftNodeIsCharacter_32(tg_io_outputs_leftNodeIsCharacter_32),
    .io_outputs_leftNodeIsCharacter_33(tg_io_outputs_leftNodeIsCharacter_33),
    .io_outputs_leftNodeIsCharacter_34(tg_io_outputs_leftNodeIsCharacter_34),
    .io_outputs_leftNodeIsCharacter_35(tg_io_outputs_leftNodeIsCharacter_35),
    .io_outputs_leftNodeIsCharacter_36(tg_io_outputs_leftNodeIsCharacter_36),
    .io_outputs_leftNodeIsCharacter_37(tg_io_outputs_leftNodeIsCharacter_37),
    .io_outputs_leftNodeIsCharacter_38(tg_io_outputs_leftNodeIsCharacter_38),
    .io_outputs_leftNodeIsCharacter_39(tg_io_outputs_leftNodeIsCharacter_39),
    .io_outputs_leftNodeIsCharacter_40(tg_io_outputs_leftNodeIsCharacter_40),
    .io_outputs_leftNodeIsCharacter_41(tg_io_outputs_leftNodeIsCharacter_41),
    .io_outputs_leftNodeIsCharacter_42(tg_io_outputs_leftNodeIsCharacter_42),
    .io_outputs_leftNodeIsCharacter_43(tg_io_outputs_leftNodeIsCharacter_43),
    .io_outputs_leftNodeIsCharacter_44(tg_io_outputs_leftNodeIsCharacter_44),
    .io_outputs_leftNodeIsCharacter_45(tg_io_outputs_leftNodeIsCharacter_45),
    .io_outputs_leftNodeIsCharacter_46(tg_io_outputs_leftNodeIsCharacter_46),
    .io_outputs_leftNodeIsCharacter_47(tg_io_outputs_leftNodeIsCharacter_47),
    .io_outputs_leftNodeIsCharacter_48(tg_io_outputs_leftNodeIsCharacter_48),
    .io_outputs_leftNodeIsCharacter_49(tg_io_outputs_leftNodeIsCharacter_49),
    .io_outputs_leftNodeIsCharacter_50(tg_io_outputs_leftNodeIsCharacter_50),
    .io_outputs_leftNodeIsCharacter_51(tg_io_outputs_leftNodeIsCharacter_51),
    .io_outputs_leftNodeIsCharacter_52(tg_io_outputs_leftNodeIsCharacter_52),
    .io_outputs_leftNodeIsCharacter_53(tg_io_outputs_leftNodeIsCharacter_53),
    .io_outputs_leftNodeIsCharacter_54(tg_io_outputs_leftNodeIsCharacter_54),
    .io_outputs_leftNodeIsCharacter_55(tg_io_outputs_leftNodeIsCharacter_55),
    .io_outputs_leftNodeIsCharacter_56(tg_io_outputs_leftNodeIsCharacter_56),
    .io_outputs_leftNodeIsCharacter_57(tg_io_outputs_leftNodeIsCharacter_57),
    .io_outputs_leftNodeIsCharacter_58(tg_io_outputs_leftNodeIsCharacter_58),
    .io_outputs_leftNodeIsCharacter_59(tg_io_outputs_leftNodeIsCharacter_59),
    .io_outputs_leftNodeIsCharacter_60(tg_io_outputs_leftNodeIsCharacter_60),
    .io_outputs_leftNodeIsCharacter_61(tg_io_outputs_leftNodeIsCharacter_61),
    .io_outputs_leftNodeIsCharacter_62(tg_io_outputs_leftNodeIsCharacter_62),
    .io_outputs_leftNodeIsCharacter_63(tg_io_outputs_leftNodeIsCharacter_63),
    .io_outputs_rightNodeIsCharacter_0(tg_io_outputs_rightNodeIsCharacter_0),
    .io_outputs_rightNodeIsCharacter_1(tg_io_outputs_rightNodeIsCharacter_1),
    .io_outputs_rightNodeIsCharacter_2(tg_io_outputs_rightNodeIsCharacter_2),
    .io_outputs_rightNodeIsCharacter_3(tg_io_outputs_rightNodeIsCharacter_3),
    .io_outputs_rightNodeIsCharacter_4(tg_io_outputs_rightNodeIsCharacter_4),
    .io_outputs_rightNodeIsCharacter_5(tg_io_outputs_rightNodeIsCharacter_5),
    .io_outputs_rightNodeIsCharacter_6(tg_io_outputs_rightNodeIsCharacter_6),
    .io_outputs_rightNodeIsCharacter_7(tg_io_outputs_rightNodeIsCharacter_7),
    .io_outputs_rightNodeIsCharacter_8(tg_io_outputs_rightNodeIsCharacter_8),
    .io_outputs_rightNodeIsCharacter_9(tg_io_outputs_rightNodeIsCharacter_9),
    .io_outputs_rightNodeIsCharacter_10(tg_io_outputs_rightNodeIsCharacter_10),
    .io_outputs_rightNodeIsCharacter_11(tg_io_outputs_rightNodeIsCharacter_11),
    .io_outputs_rightNodeIsCharacter_12(tg_io_outputs_rightNodeIsCharacter_12),
    .io_outputs_rightNodeIsCharacter_13(tg_io_outputs_rightNodeIsCharacter_13),
    .io_outputs_rightNodeIsCharacter_14(tg_io_outputs_rightNodeIsCharacter_14),
    .io_outputs_rightNodeIsCharacter_15(tg_io_outputs_rightNodeIsCharacter_15),
    .io_outputs_rightNodeIsCharacter_16(tg_io_outputs_rightNodeIsCharacter_16),
    .io_outputs_rightNodeIsCharacter_17(tg_io_outputs_rightNodeIsCharacter_17),
    .io_outputs_rightNodeIsCharacter_18(tg_io_outputs_rightNodeIsCharacter_18),
    .io_outputs_rightNodeIsCharacter_19(tg_io_outputs_rightNodeIsCharacter_19),
    .io_outputs_rightNodeIsCharacter_20(tg_io_outputs_rightNodeIsCharacter_20),
    .io_outputs_rightNodeIsCharacter_21(tg_io_outputs_rightNodeIsCharacter_21),
    .io_outputs_rightNodeIsCharacter_22(tg_io_outputs_rightNodeIsCharacter_22),
    .io_outputs_rightNodeIsCharacter_23(tg_io_outputs_rightNodeIsCharacter_23),
    .io_outputs_rightNodeIsCharacter_24(tg_io_outputs_rightNodeIsCharacter_24),
    .io_outputs_rightNodeIsCharacter_25(tg_io_outputs_rightNodeIsCharacter_25),
    .io_outputs_rightNodeIsCharacter_26(tg_io_outputs_rightNodeIsCharacter_26),
    .io_outputs_rightNodeIsCharacter_27(tg_io_outputs_rightNodeIsCharacter_27),
    .io_outputs_rightNodeIsCharacter_28(tg_io_outputs_rightNodeIsCharacter_28),
    .io_outputs_rightNodeIsCharacter_29(tg_io_outputs_rightNodeIsCharacter_29),
    .io_outputs_rightNodeIsCharacter_30(tg_io_outputs_rightNodeIsCharacter_30),
    .io_outputs_rightNodeIsCharacter_31(tg_io_outputs_rightNodeIsCharacter_31),
    .io_outputs_rightNodeIsCharacter_32(tg_io_outputs_rightNodeIsCharacter_32),
    .io_outputs_rightNodeIsCharacter_33(tg_io_outputs_rightNodeIsCharacter_33),
    .io_outputs_rightNodeIsCharacter_34(tg_io_outputs_rightNodeIsCharacter_34),
    .io_outputs_rightNodeIsCharacter_35(tg_io_outputs_rightNodeIsCharacter_35),
    .io_outputs_rightNodeIsCharacter_36(tg_io_outputs_rightNodeIsCharacter_36),
    .io_outputs_rightNodeIsCharacter_37(tg_io_outputs_rightNodeIsCharacter_37),
    .io_outputs_rightNodeIsCharacter_38(tg_io_outputs_rightNodeIsCharacter_38),
    .io_outputs_rightNodeIsCharacter_39(tg_io_outputs_rightNodeIsCharacter_39),
    .io_outputs_rightNodeIsCharacter_40(tg_io_outputs_rightNodeIsCharacter_40),
    .io_outputs_rightNodeIsCharacter_41(tg_io_outputs_rightNodeIsCharacter_41),
    .io_outputs_rightNodeIsCharacter_42(tg_io_outputs_rightNodeIsCharacter_42),
    .io_outputs_rightNodeIsCharacter_43(tg_io_outputs_rightNodeIsCharacter_43),
    .io_outputs_rightNodeIsCharacter_44(tg_io_outputs_rightNodeIsCharacter_44),
    .io_outputs_rightNodeIsCharacter_45(tg_io_outputs_rightNodeIsCharacter_45),
    .io_outputs_rightNodeIsCharacter_46(tg_io_outputs_rightNodeIsCharacter_46),
    .io_outputs_rightNodeIsCharacter_47(tg_io_outputs_rightNodeIsCharacter_47),
    .io_outputs_rightNodeIsCharacter_48(tg_io_outputs_rightNodeIsCharacter_48),
    .io_outputs_rightNodeIsCharacter_49(tg_io_outputs_rightNodeIsCharacter_49),
    .io_outputs_rightNodeIsCharacter_50(tg_io_outputs_rightNodeIsCharacter_50),
    .io_outputs_rightNodeIsCharacter_51(tg_io_outputs_rightNodeIsCharacter_51),
    .io_outputs_rightNodeIsCharacter_52(tg_io_outputs_rightNodeIsCharacter_52),
    .io_outputs_rightNodeIsCharacter_53(tg_io_outputs_rightNodeIsCharacter_53),
    .io_outputs_rightNodeIsCharacter_54(tg_io_outputs_rightNodeIsCharacter_54),
    .io_outputs_rightNodeIsCharacter_55(tg_io_outputs_rightNodeIsCharacter_55),
    .io_outputs_rightNodeIsCharacter_56(tg_io_outputs_rightNodeIsCharacter_56),
    .io_outputs_rightNodeIsCharacter_57(tg_io_outputs_rightNodeIsCharacter_57),
    .io_outputs_rightNodeIsCharacter_58(tg_io_outputs_rightNodeIsCharacter_58),
    .io_outputs_rightNodeIsCharacter_59(tg_io_outputs_rightNodeIsCharacter_59),
    .io_outputs_rightNodeIsCharacter_60(tg_io_outputs_rightNodeIsCharacter_60),
    .io_outputs_rightNodeIsCharacter_61(tg_io_outputs_rightNodeIsCharacter_61),
    .io_outputs_rightNodeIsCharacter_62(tg_io_outputs_rightNodeIsCharacter_62),
    .io_outputs_rightNodeIsCharacter_63(tg_io_outputs_rightNodeIsCharacter_63),
    .io_outputs_validNodes(tg_io_outputs_validNodes),
    .io_outputs_validCharacters(tg_io_outputs_validCharacters),
    .io_finished(tg_io_finished)
  );
  treeDepthCounter tdc ( // @[topLevel.scala 57:19]
    .clock(tdc_clock),
    .reset(tdc_reset),
    .io_start(tdc_io_start),
    .io_inputs_leftNode_0(tdc_io_inputs_leftNode_0),
    .io_inputs_leftNode_1(tdc_io_inputs_leftNode_1),
    .io_inputs_leftNode_2(tdc_io_inputs_leftNode_2),
    .io_inputs_leftNode_3(tdc_io_inputs_leftNode_3),
    .io_inputs_leftNode_4(tdc_io_inputs_leftNode_4),
    .io_inputs_leftNode_5(tdc_io_inputs_leftNode_5),
    .io_inputs_leftNode_6(tdc_io_inputs_leftNode_6),
    .io_inputs_leftNode_7(tdc_io_inputs_leftNode_7),
    .io_inputs_leftNode_8(tdc_io_inputs_leftNode_8),
    .io_inputs_leftNode_9(tdc_io_inputs_leftNode_9),
    .io_inputs_leftNode_10(tdc_io_inputs_leftNode_10),
    .io_inputs_leftNode_11(tdc_io_inputs_leftNode_11),
    .io_inputs_leftNode_12(tdc_io_inputs_leftNode_12),
    .io_inputs_leftNode_13(tdc_io_inputs_leftNode_13),
    .io_inputs_leftNode_14(tdc_io_inputs_leftNode_14),
    .io_inputs_leftNode_15(tdc_io_inputs_leftNode_15),
    .io_inputs_leftNode_16(tdc_io_inputs_leftNode_16),
    .io_inputs_leftNode_17(tdc_io_inputs_leftNode_17),
    .io_inputs_leftNode_18(tdc_io_inputs_leftNode_18),
    .io_inputs_leftNode_19(tdc_io_inputs_leftNode_19),
    .io_inputs_leftNode_20(tdc_io_inputs_leftNode_20),
    .io_inputs_leftNode_21(tdc_io_inputs_leftNode_21),
    .io_inputs_leftNode_22(tdc_io_inputs_leftNode_22),
    .io_inputs_leftNode_23(tdc_io_inputs_leftNode_23),
    .io_inputs_leftNode_24(tdc_io_inputs_leftNode_24),
    .io_inputs_leftNode_25(tdc_io_inputs_leftNode_25),
    .io_inputs_leftNode_26(tdc_io_inputs_leftNode_26),
    .io_inputs_leftNode_27(tdc_io_inputs_leftNode_27),
    .io_inputs_leftNode_28(tdc_io_inputs_leftNode_28),
    .io_inputs_leftNode_29(tdc_io_inputs_leftNode_29),
    .io_inputs_leftNode_30(tdc_io_inputs_leftNode_30),
    .io_inputs_leftNode_31(tdc_io_inputs_leftNode_31),
    .io_inputs_leftNode_32(tdc_io_inputs_leftNode_32),
    .io_inputs_leftNode_33(tdc_io_inputs_leftNode_33),
    .io_inputs_leftNode_34(tdc_io_inputs_leftNode_34),
    .io_inputs_leftNode_35(tdc_io_inputs_leftNode_35),
    .io_inputs_leftNode_36(tdc_io_inputs_leftNode_36),
    .io_inputs_leftNode_37(tdc_io_inputs_leftNode_37),
    .io_inputs_leftNode_38(tdc_io_inputs_leftNode_38),
    .io_inputs_leftNode_39(tdc_io_inputs_leftNode_39),
    .io_inputs_leftNode_40(tdc_io_inputs_leftNode_40),
    .io_inputs_leftNode_41(tdc_io_inputs_leftNode_41),
    .io_inputs_leftNode_42(tdc_io_inputs_leftNode_42),
    .io_inputs_leftNode_43(tdc_io_inputs_leftNode_43),
    .io_inputs_leftNode_44(tdc_io_inputs_leftNode_44),
    .io_inputs_leftNode_45(tdc_io_inputs_leftNode_45),
    .io_inputs_leftNode_46(tdc_io_inputs_leftNode_46),
    .io_inputs_leftNode_47(tdc_io_inputs_leftNode_47),
    .io_inputs_leftNode_48(tdc_io_inputs_leftNode_48),
    .io_inputs_leftNode_49(tdc_io_inputs_leftNode_49),
    .io_inputs_leftNode_50(tdc_io_inputs_leftNode_50),
    .io_inputs_leftNode_51(tdc_io_inputs_leftNode_51),
    .io_inputs_leftNode_52(tdc_io_inputs_leftNode_52),
    .io_inputs_leftNode_53(tdc_io_inputs_leftNode_53),
    .io_inputs_leftNode_54(tdc_io_inputs_leftNode_54),
    .io_inputs_leftNode_55(tdc_io_inputs_leftNode_55),
    .io_inputs_leftNode_56(tdc_io_inputs_leftNode_56),
    .io_inputs_leftNode_57(tdc_io_inputs_leftNode_57),
    .io_inputs_leftNode_58(tdc_io_inputs_leftNode_58),
    .io_inputs_leftNode_59(tdc_io_inputs_leftNode_59),
    .io_inputs_leftNode_60(tdc_io_inputs_leftNode_60),
    .io_inputs_leftNode_61(tdc_io_inputs_leftNode_61),
    .io_inputs_leftNode_62(tdc_io_inputs_leftNode_62),
    .io_inputs_leftNode_63(tdc_io_inputs_leftNode_63),
    .io_inputs_rightNode_0(tdc_io_inputs_rightNode_0),
    .io_inputs_rightNode_1(tdc_io_inputs_rightNode_1),
    .io_inputs_rightNode_2(tdc_io_inputs_rightNode_2),
    .io_inputs_rightNode_3(tdc_io_inputs_rightNode_3),
    .io_inputs_rightNode_4(tdc_io_inputs_rightNode_4),
    .io_inputs_rightNode_5(tdc_io_inputs_rightNode_5),
    .io_inputs_rightNode_6(tdc_io_inputs_rightNode_6),
    .io_inputs_rightNode_7(tdc_io_inputs_rightNode_7),
    .io_inputs_rightNode_8(tdc_io_inputs_rightNode_8),
    .io_inputs_rightNode_9(tdc_io_inputs_rightNode_9),
    .io_inputs_rightNode_10(tdc_io_inputs_rightNode_10),
    .io_inputs_rightNode_11(tdc_io_inputs_rightNode_11),
    .io_inputs_rightNode_12(tdc_io_inputs_rightNode_12),
    .io_inputs_rightNode_13(tdc_io_inputs_rightNode_13),
    .io_inputs_rightNode_14(tdc_io_inputs_rightNode_14),
    .io_inputs_rightNode_15(tdc_io_inputs_rightNode_15),
    .io_inputs_rightNode_16(tdc_io_inputs_rightNode_16),
    .io_inputs_rightNode_17(tdc_io_inputs_rightNode_17),
    .io_inputs_rightNode_18(tdc_io_inputs_rightNode_18),
    .io_inputs_rightNode_19(tdc_io_inputs_rightNode_19),
    .io_inputs_rightNode_20(tdc_io_inputs_rightNode_20),
    .io_inputs_rightNode_21(tdc_io_inputs_rightNode_21),
    .io_inputs_rightNode_22(tdc_io_inputs_rightNode_22),
    .io_inputs_rightNode_23(tdc_io_inputs_rightNode_23),
    .io_inputs_rightNode_24(tdc_io_inputs_rightNode_24),
    .io_inputs_rightNode_25(tdc_io_inputs_rightNode_25),
    .io_inputs_rightNode_26(tdc_io_inputs_rightNode_26),
    .io_inputs_rightNode_27(tdc_io_inputs_rightNode_27),
    .io_inputs_rightNode_28(tdc_io_inputs_rightNode_28),
    .io_inputs_rightNode_29(tdc_io_inputs_rightNode_29),
    .io_inputs_rightNode_30(tdc_io_inputs_rightNode_30),
    .io_inputs_rightNode_31(tdc_io_inputs_rightNode_31),
    .io_inputs_rightNode_32(tdc_io_inputs_rightNode_32),
    .io_inputs_rightNode_33(tdc_io_inputs_rightNode_33),
    .io_inputs_rightNode_34(tdc_io_inputs_rightNode_34),
    .io_inputs_rightNode_35(tdc_io_inputs_rightNode_35),
    .io_inputs_rightNode_36(tdc_io_inputs_rightNode_36),
    .io_inputs_rightNode_37(tdc_io_inputs_rightNode_37),
    .io_inputs_rightNode_38(tdc_io_inputs_rightNode_38),
    .io_inputs_rightNode_39(tdc_io_inputs_rightNode_39),
    .io_inputs_rightNode_40(tdc_io_inputs_rightNode_40),
    .io_inputs_rightNode_41(tdc_io_inputs_rightNode_41),
    .io_inputs_rightNode_42(tdc_io_inputs_rightNode_42),
    .io_inputs_rightNode_43(tdc_io_inputs_rightNode_43),
    .io_inputs_rightNode_44(tdc_io_inputs_rightNode_44),
    .io_inputs_rightNode_45(tdc_io_inputs_rightNode_45),
    .io_inputs_rightNode_46(tdc_io_inputs_rightNode_46),
    .io_inputs_rightNode_47(tdc_io_inputs_rightNode_47),
    .io_inputs_rightNode_48(tdc_io_inputs_rightNode_48),
    .io_inputs_rightNode_49(tdc_io_inputs_rightNode_49),
    .io_inputs_rightNode_50(tdc_io_inputs_rightNode_50),
    .io_inputs_rightNode_51(tdc_io_inputs_rightNode_51),
    .io_inputs_rightNode_52(tdc_io_inputs_rightNode_52),
    .io_inputs_rightNode_53(tdc_io_inputs_rightNode_53),
    .io_inputs_rightNode_54(tdc_io_inputs_rightNode_54),
    .io_inputs_rightNode_55(tdc_io_inputs_rightNode_55),
    .io_inputs_rightNode_56(tdc_io_inputs_rightNode_56),
    .io_inputs_rightNode_57(tdc_io_inputs_rightNode_57),
    .io_inputs_rightNode_58(tdc_io_inputs_rightNode_58),
    .io_inputs_rightNode_59(tdc_io_inputs_rightNode_59),
    .io_inputs_rightNode_60(tdc_io_inputs_rightNode_60),
    .io_inputs_rightNode_61(tdc_io_inputs_rightNode_61),
    .io_inputs_rightNode_62(tdc_io_inputs_rightNode_62),
    .io_inputs_rightNode_63(tdc_io_inputs_rightNode_63),
    .io_inputs_leftNodeIsCharacter_0(tdc_io_inputs_leftNodeIsCharacter_0),
    .io_inputs_leftNodeIsCharacter_1(tdc_io_inputs_leftNodeIsCharacter_1),
    .io_inputs_leftNodeIsCharacter_2(tdc_io_inputs_leftNodeIsCharacter_2),
    .io_inputs_leftNodeIsCharacter_3(tdc_io_inputs_leftNodeIsCharacter_3),
    .io_inputs_leftNodeIsCharacter_4(tdc_io_inputs_leftNodeIsCharacter_4),
    .io_inputs_leftNodeIsCharacter_5(tdc_io_inputs_leftNodeIsCharacter_5),
    .io_inputs_leftNodeIsCharacter_6(tdc_io_inputs_leftNodeIsCharacter_6),
    .io_inputs_leftNodeIsCharacter_7(tdc_io_inputs_leftNodeIsCharacter_7),
    .io_inputs_leftNodeIsCharacter_8(tdc_io_inputs_leftNodeIsCharacter_8),
    .io_inputs_leftNodeIsCharacter_9(tdc_io_inputs_leftNodeIsCharacter_9),
    .io_inputs_leftNodeIsCharacter_10(tdc_io_inputs_leftNodeIsCharacter_10),
    .io_inputs_leftNodeIsCharacter_11(tdc_io_inputs_leftNodeIsCharacter_11),
    .io_inputs_leftNodeIsCharacter_12(tdc_io_inputs_leftNodeIsCharacter_12),
    .io_inputs_leftNodeIsCharacter_13(tdc_io_inputs_leftNodeIsCharacter_13),
    .io_inputs_leftNodeIsCharacter_14(tdc_io_inputs_leftNodeIsCharacter_14),
    .io_inputs_leftNodeIsCharacter_15(tdc_io_inputs_leftNodeIsCharacter_15),
    .io_inputs_leftNodeIsCharacter_16(tdc_io_inputs_leftNodeIsCharacter_16),
    .io_inputs_leftNodeIsCharacter_17(tdc_io_inputs_leftNodeIsCharacter_17),
    .io_inputs_leftNodeIsCharacter_18(tdc_io_inputs_leftNodeIsCharacter_18),
    .io_inputs_leftNodeIsCharacter_19(tdc_io_inputs_leftNodeIsCharacter_19),
    .io_inputs_leftNodeIsCharacter_20(tdc_io_inputs_leftNodeIsCharacter_20),
    .io_inputs_leftNodeIsCharacter_21(tdc_io_inputs_leftNodeIsCharacter_21),
    .io_inputs_leftNodeIsCharacter_22(tdc_io_inputs_leftNodeIsCharacter_22),
    .io_inputs_leftNodeIsCharacter_23(tdc_io_inputs_leftNodeIsCharacter_23),
    .io_inputs_leftNodeIsCharacter_24(tdc_io_inputs_leftNodeIsCharacter_24),
    .io_inputs_leftNodeIsCharacter_25(tdc_io_inputs_leftNodeIsCharacter_25),
    .io_inputs_leftNodeIsCharacter_26(tdc_io_inputs_leftNodeIsCharacter_26),
    .io_inputs_leftNodeIsCharacter_27(tdc_io_inputs_leftNodeIsCharacter_27),
    .io_inputs_leftNodeIsCharacter_28(tdc_io_inputs_leftNodeIsCharacter_28),
    .io_inputs_leftNodeIsCharacter_29(tdc_io_inputs_leftNodeIsCharacter_29),
    .io_inputs_leftNodeIsCharacter_30(tdc_io_inputs_leftNodeIsCharacter_30),
    .io_inputs_leftNodeIsCharacter_31(tdc_io_inputs_leftNodeIsCharacter_31),
    .io_inputs_leftNodeIsCharacter_32(tdc_io_inputs_leftNodeIsCharacter_32),
    .io_inputs_leftNodeIsCharacter_33(tdc_io_inputs_leftNodeIsCharacter_33),
    .io_inputs_leftNodeIsCharacter_34(tdc_io_inputs_leftNodeIsCharacter_34),
    .io_inputs_leftNodeIsCharacter_35(tdc_io_inputs_leftNodeIsCharacter_35),
    .io_inputs_leftNodeIsCharacter_36(tdc_io_inputs_leftNodeIsCharacter_36),
    .io_inputs_leftNodeIsCharacter_37(tdc_io_inputs_leftNodeIsCharacter_37),
    .io_inputs_leftNodeIsCharacter_38(tdc_io_inputs_leftNodeIsCharacter_38),
    .io_inputs_leftNodeIsCharacter_39(tdc_io_inputs_leftNodeIsCharacter_39),
    .io_inputs_leftNodeIsCharacter_40(tdc_io_inputs_leftNodeIsCharacter_40),
    .io_inputs_leftNodeIsCharacter_41(tdc_io_inputs_leftNodeIsCharacter_41),
    .io_inputs_leftNodeIsCharacter_42(tdc_io_inputs_leftNodeIsCharacter_42),
    .io_inputs_leftNodeIsCharacter_43(tdc_io_inputs_leftNodeIsCharacter_43),
    .io_inputs_leftNodeIsCharacter_44(tdc_io_inputs_leftNodeIsCharacter_44),
    .io_inputs_leftNodeIsCharacter_45(tdc_io_inputs_leftNodeIsCharacter_45),
    .io_inputs_leftNodeIsCharacter_46(tdc_io_inputs_leftNodeIsCharacter_46),
    .io_inputs_leftNodeIsCharacter_47(tdc_io_inputs_leftNodeIsCharacter_47),
    .io_inputs_leftNodeIsCharacter_48(tdc_io_inputs_leftNodeIsCharacter_48),
    .io_inputs_leftNodeIsCharacter_49(tdc_io_inputs_leftNodeIsCharacter_49),
    .io_inputs_leftNodeIsCharacter_50(tdc_io_inputs_leftNodeIsCharacter_50),
    .io_inputs_leftNodeIsCharacter_51(tdc_io_inputs_leftNodeIsCharacter_51),
    .io_inputs_leftNodeIsCharacter_52(tdc_io_inputs_leftNodeIsCharacter_52),
    .io_inputs_leftNodeIsCharacter_53(tdc_io_inputs_leftNodeIsCharacter_53),
    .io_inputs_leftNodeIsCharacter_54(tdc_io_inputs_leftNodeIsCharacter_54),
    .io_inputs_leftNodeIsCharacter_55(tdc_io_inputs_leftNodeIsCharacter_55),
    .io_inputs_leftNodeIsCharacter_56(tdc_io_inputs_leftNodeIsCharacter_56),
    .io_inputs_leftNodeIsCharacter_57(tdc_io_inputs_leftNodeIsCharacter_57),
    .io_inputs_leftNodeIsCharacter_58(tdc_io_inputs_leftNodeIsCharacter_58),
    .io_inputs_leftNodeIsCharacter_59(tdc_io_inputs_leftNodeIsCharacter_59),
    .io_inputs_leftNodeIsCharacter_60(tdc_io_inputs_leftNodeIsCharacter_60),
    .io_inputs_leftNodeIsCharacter_61(tdc_io_inputs_leftNodeIsCharacter_61),
    .io_inputs_leftNodeIsCharacter_62(tdc_io_inputs_leftNodeIsCharacter_62),
    .io_inputs_leftNodeIsCharacter_63(tdc_io_inputs_leftNodeIsCharacter_63),
    .io_inputs_rightNodeIsCharacter_0(tdc_io_inputs_rightNodeIsCharacter_0),
    .io_inputs_rightNodeIsCharacter_1(tdc_io_inputs_rightNodeIsCharacter_1),
    .io_inputs_rightNodeIsCharacter_2(tdc_io_inputs_rightNodeIsCharacter_2),
    .io_inputs_rightNodeIsCharacter_3(tdc_io_inputs_rightNodeIsCharacter_3),
    .io_inputs_rightNodeIsCharacter_4(tdc_io_inputs_rightNodeIsCharacter_4),
    .io_inputs_rightNodeIsCharacter_5(tdc_io_inputs_rightNodeIsCharacter_5),
    .io_inputs_rightNodeIsCharacter_6(tdc_io_inputs_rightNodeIsCharacter_6),
    .io_inputs_rightNodeIsCharacter_7(tdc_io_inputs_rightNodeIsCharacter_7),
    .io_inputs_rightNodeIsCharacter_8(tdc_io_inputs_rightNodeIsCharacter_8),
    .io_inputs_rightNodeIsCharacter_9(tdc_io_inputs_rightNodeIsCharacter_9),
    .io_inputs_rightNodeIsCharacter_10(tdc_io_inputs_rightNodeIsCharacter_10),
    .io_inputs_rightNodeIsCharacter_11(tdc_io_inputs_rightNodeIsCharacter_11),
    .io_inputs_rightNodeIsCharacter_12(tdc_io_inputs_rightNodeIsCharacter_12),
    .io_inputs_rightNodeIsCharacter_13(tdc_io_inputs_rightNodeIsCharacter_13),
    .io_inputs_rightNodeIsCharacter_14(tdc_io_inputs_rightNodeIsCharacter_14),
    .io_inputs_rightNodeIsCharacter_15(tdc_io_inputs_rightNodeIsCharacter_15),
    .io_inputs_rightNodeIsCharacter_16(tdc_io_inputs_rightNodeIsCharacter_16),
    .io_inputs_rightNodeIsCharacter_17(tdc_io_inputs_rightNodeIsCharacter_17),
    .io_inputs_rightNodeIsCharacter_18(tdc_io_inputs_rightNodeIsCharacter_18),
    .io_inputs_rightNodeIsCharacter_19(tdc_io_inputs_rightNodeIsCharacter_19),
    .io_inputs_rightNodeIsCharacter_20(tdc_io_inputs_rightNodeIsCharacter_20),
    .io_inputs_rightNodeIsCharacter_21(tdc_io_inputs_rightNodeIsCharacter_21),
    .io_inputs_rightNodeIsCharacter_22(tdc_io_inputs_rightNodeIsCharacter_22),
    .io_inputs_rightNodeIsCharacter_23(tdc_io_inputs_rightNodeIsCharacter_23),
    .io_inputs_rightNodeIsCharacter_24(tdc_io_inputs_rightNodeIsCharacter_24),
    .io_inputs_rightNodeIsCharacter_25(tdc_io_inputs_rightNodeIsCharacter_25),
    .io_inputs_rightNodeIsCharacter_26(tdc_io_inputs_rightNodeIsCharacter_26),
    .io_inputs_rightNodeIsCharacter_27(tdc_io_inputs_rightNodeIsCharacter_27),
    .io_inputs_rightNodeIsCharacter_28(tdc_io_inputs_rightNodeIsCharacter_28),
    .io_inputs_rightNodeIsCharacter_29(tdc_io_inputs_rightNodeIsCharacter_29),
    .io_inputs_rightNodeIsCharacter_30(tdc_io_inputs_rightNodeIsCharacter_30),
    .io_inputs_rightNodeIsCharacter_31(tdc_io_inputs_rightNodeIsCharacter_31),
    .io_inputs_rightNodeIsCharacter_32(tdc_io_inputs_rightNodeIsCharacter_32),
    .io_inputs_rightNodeIsCharacter_33(tdc_io_inputs_rightNodeIsCharacter_33),
    .io_inputs_rightNodeIsCharacter_34(tdc_io_inputs_rightNodeIsCharacter_34),
    .io_inputs_rightNodeIsCharacter_35(tdc_io_inputs_rightNodeIsCharacter_35),
    .io_inputs_rightNodeIsCharacter_36(tdc_io_inputs_rightNodeIsCharacter_36),
    .io_inputs_rightNodeIsCharacter_37(tdc_io_inputs_rightNodeIsCharacter_37),
    .io_inputs_rightNodeIsCharacter_38(tdc_io_inputs_rightNodeIsCharacter_38),
    .io_inputs_rightNodeIsCharacter_39(tdc_io_inputs_rightNodeIsCharacter_39),
    .io_inputs_rightNodeIsCharacter_40(tdc_io_inputs_rightNodeIsCharacter_40),
    .io_inputs_rightNodeIsCharacter_41(tdc_io_inputs_rightNodeIsCharacter_41),
    .io_inputs_rightNodeIsCharacter_42(tdc_io_inputs_rightNodeIsCharacter_42),
    .io_inputs_rightNodeIsCharacter_43(tdc_io_inputs_rightNodeIsCharacter_43),
    .io_inputs_rightNodeIsCharacter_44(tdc_io_inputs_rightNodeIsCharacter_44),
    .io_inputs_rightNodeIsCharacter_45(tdc_io_inputs_rightNodeIsCharacter_45),
    .io_inputs_rightNodeIsCharacter_46(tdc_io_inputs_rightNodeIsCharacter_46),
    .io_inputs_rightNodeIsCharacter_47(tdc_io_inputs_rightNodeIsCharacter_47),
    .io_inputs_rightNodeIsCharacter_48(tdc_io_inputs_rightNodeIsCharacter_48),
    .io_inputs_rightNodeIsCharacter_49(tdc_io_inputs_rightNodeIsCharacter_49),
    .io_inputs_rightNodeIsCharacter_50(tdc_io_inputs_rightNodeIsCharacter_50),
    .io_inputs_rightNodeIsCharacter_51(tdc_io_inputs_rightNodeIsCharacter_51),
    .io_inputs_rightNodeIsCharacter_52(tdc_io_inputs_rightNodeIsCharacter_52),
    .io_inputs_rightNodeIsCharacter_53(tdc_io_inputs_rightNodeIsCharacter_53),
    .io_inputs_rightNodeIsCharacter_54(tdc_io_inputs_rightNodeIsCharacter_54),
    .io_inputs_rightNodeIsCharacter_55(tdc_io_inputs_rightNodeIsCharacter_55),
    .io_inputs_rightNodeIsCharacter_56(tdc_io_inputs_rightNodeIsCharacter_56),
    .io_inputs_rightNodeIsCharacter_57(tdc_io_inputs_rightNodeIsCharacter_57),
    .io_inputs_rightNodeIsCharacter_58(tdc_io_inputs_rightNodeIsCharacter_58),
    .io_inputs_rightNodeIsCharacter_59(tdc_io_inputs_rightNodeIsCharacter_59),
    .io_inputs_rightNodeIsCharacter_60(tdc_io_inputs_rightNodeIsCharacter_60),
    .io_inputs_rightNodeIsCharacter_61(tdc_io_inputs_rightNodeIsCharacter_61),
    .io_inputs_rightNodeIsCharacter_62(tdc_io_inputs_rightNodeIsCharacter_62),
    .io_inputs_rightNodeIsCharacter_63(tdc_io_inputs_rightNodeIsCharacter_63),
    .io_inputs_validNodes(tdc_io_inputs_validNodes),
    .io_inputs_validCharacters(tdc_io_inputs_validCharacters),
    .io_outputs_characters_0(tdc_io_outputs_characters_0),
    .io_outputs_characters_1(tdc_io_outputs_characters_1),
    .io_outputs_characters_2(tdc_io_outputs_characters_2),
    .io_outputs_characters_3(tdc_io_outputs_characters_3),
    .io_outputs_characters_4(tdc_io_outputs_characters_4),
    .io_outputs_characters_5(tdc_io_outputs_characters_5),
    .io_outputs_characters_6(tdc_io_outputs_characters_6),
    .io_outputs_characters_7(tdc_io_outputs_characters_7),
    .io_outputs_characters_8(tdc_io_outputs_characters_8),
    .io_outputs_characters_9(tdc_io_outputs_characters_9),
    .io_outputs_characters_10(tdc_io_outputs_characters_10),
    .io_outputs_characters_11(tdc_io_outputs_characters_11),
    .io_outputs_characters_12(tdc_io_outputs_characters_12),
    .io_outputs_characters_13(tdc_io_outputs_characters_13),
    .io_outputs_characters_14(tdc_io_outputs_characters_14),
    .io_outputs_characters_15(tdc_io_outputs_characters_15),
    .io_outputs_characters_16(tdc_io_outputs_characters_16),
    .io_outputs_characters_17(tdc_io_outputs_characters_17),
    .io_outputs_characters_18(tdc_io_outputs_characters_18),
    .io_outputs_characters_19(tdc_io_outputs_characters_19),
    .io_outputs_characters_20(tdc_io_outputs_characters_20),
    .io_outputs_characters_21(tdc_io_outputs_characters_21),
    .io_outputs_characters_22(tdc_io_outputs_characters_22),
    .io_outputs_characters_23(tdc_io_outputs_characters_23),
    .io_outputs_characters_24(tdc_io_outputs_characters_24),
    .io_outputs_characters_25(tdc_io_outputs_characters_25),
    .io_outputs_characters_26(tdc_io_outputs_characters_26),
    .io_outputs_characters_27(tdc_io_outputs_characters_27),
    .io_outputs_characters_28(tdc_io_outputs_characters_28),
    .io_outputs_characters_29(tdc_io_outputs_characters_29),
    .io_outputs_characters_30(tdc_io_outputs_characters_30),
    .io_outputs_characters_31(tdc_io_outputs_characters_31),
    .io_outputs_depths_0(tdc_io_outputs_depths_0),
    .io_outputs_depths_1(tdc_io_outputs_depths_1),
    .io_outputs_depths_2(tdc_io_outputs_depths_2),
    .io_outputs_depths_3(tdc_io_outputs_depths_3),
    .io_outputs_depths_4(tdc_io_outputs_depths_4),
    .io_outputs_depths_5(tdc_io_outputs_depths_5),
    .io_outputs_depths_6(tdc_io_outputs_depths_6),
    .io_outputs_depths_7(tdc_io_outputs_depths_7),
    .io_outputs_depths_8(tdc_io_outputs_depths_8),
    .io_outputs_depths_9(tdc_io_outputs_depths_9),
    .io_outputs_depths_10(tdc_io_outputs_depths_10),
    .io_outputs_depths_11(tdc_io_outputs_depths_11),
    .io_outputs_depths_12(tdc_io_outputs_depths_12),
    .io_outputs_depths_13(tdc_io_outputs_depths_13),
    .io_outputs_depths_14(tdc_io_outputs_depths_14),
    .io_outputs_depths_15(tdc_io_outputs_depths_15),
    .io_outputs_depths_16(tdc_io_outputs_depths_16),
    .io_outputs_depths_17(tdc_io_outputs_depths_17),
    .io_outputs_depths_18(tdc_io_outputs_depths_18),
    .io_outputs_depths_19(tdc_io_outputs_depths_19),
    .io_outputs_depths_20(tdc_io_outputs_depths_20),
    .io_outputs_depths_21(tdc_io_outputs_depths_21),
    .io_outputs_depths_22(tdc_io_outputs_depths_22),
    .io_outputs_depths_23(tdc_io_outputs_depths_23),
    .io_outputs_depths_24(tdc_io_outputs_depths_24),
    .io_outputs_depths_25(tdc_io_outputs_depths_25),
    .io_outputs_depths_26(tdc_io_outputs_depths_26),
    .io_outputs_depths_27(tdc_io_outputs_depths_27),
    .io_outputs_depths_28(tdc_io_outputs_depths_28),
    .io_outputs_depths_29(tdc_io_outputs_depths_29),
    .io_outputs_depths_30(tdc_io_outputs_depths_30),
    .io_outputs_depths_31(tdc_io_outputs_depths_31),
    .io_outputs_validCharacters(tdc_io_outputs_validCharacters),
    .io_finished(tdc_io_finished)
  );
  sort sltg ( // @[topLevel.scala 58:20]
    .clock(sltg_clock),
    .reset(sltg_reset),
    .io_start(sltg_io_start),
    .io_inputs_characters_0(sltg_io_inputs_characters_0),
    .io_inputs_characters_1(sltg_io_inputs_characters_1),
    .io_inputs_characters_2(sltg_io_inputs_characters_2),
    .io_inputs_characters_3(sltg_io_inputs_characters_3),
    .io_inputs_characters_4(sltg_io_inputs_characters_4),
    .io_inputs_characters_5(sltg_io_inputs_characters_5),
    .io_inputs_characters_6(sltg_io_inputs_characters_6),
    .io_inputs_characters_7(sltg_io_inputs_characters_7),
    .io_inputs_characters_8(sltg_io_inputs_characters_8),
    .io_inputs_characters_9(sltg_io_inputs_characters_9),
    .io_inputs_characters_10(sltg_io_inputs_characters_10),
    .io_inputs_characters_11(sltg_io_inputs_characters_11),
    .io_inputs_characters_12(sltg_io_inputs_characters_12),
    .io_inputs_characters_13(sltg_io_inputs_characters_13),
    .io_inputs_characters_14(sltg_io_inputs_characters_14),
    .io_inputs_characters_15(sltg_io_inputs_characters_15),
    .io_inputs_characters_16(sltg_io_inputs_characters_16),
    .io_inputs_characters_17(sltg_io_inputs_characters_17),
    .io_inputs_characters_18(sltg_io_inputs_characters_18),
    .io_inputs_characters_19(sltg_io_inputs_characters_19),
    .io_inputs_characters_20(sltg_io_inputs_characters_20),
    .io_inputs_characters_21(sltg_io_inputs_characters_21),
    .io_inputs_characters_22(sltg_io_inputs_characters_22),
    .io_inputs_characters_23(sltg_io_inputs_characters_23),
    .io_inputs_characters_24(sltg_io_inputs_characters_24),
    .io_inputs_characters_25(sltg_io_inputs_characters_25),
    .io_inputs_characters_26(sltg_io_inputs_characters_26),
    .io_inputs_characters_27(sltg_io_inputs_characters_27),
    .io_inputs_characters_28(sltg_io_inputs_characters_28),
    .io_inputs_characters_29(sltg_io_inputs_characters_29),
    .io_inputs_characters_30(sltg_io_inputs_characters_30),
    .io_inputs_characters_31(sltg_io_inputs_characters_31),
    .io_inputs_depths_0(sltg_io_inputs_depths_0),
    .io_inputs_depths_1(sltg_io_inputs_depths_1),
    .io_inputs_depths_2(sltg_io_inputs_depths_2),
    .io_inputs_depths_3(sltg_io_inputs_depths_3),
    .io_inputs_depths_4(sltg_io_inputs_depths_4),
    .io_inputs_depths_5(sltg_io_inputs_depths_5),
    .io_inputs_depths_6(sltg_io_inputs_depths_6),
    .io_inputs_depths_7(sltg_io_inputs_depths_7),
    .io_inputs_depths_8(sltg_io_inputs_depths_8),
    .io_inputs_depths_9(sltg_io_inputs_depths_9),
    .io_inputs_depths_10(sltg_io_inputs_depths_10),
    .io_inputs_depths_11(sltg_io_inputs_depths_11),
    .io_inputs_depths_12(sltg_io_inputs_depths_12),
    .io_inputs_depths_13(sltg_io_inputs_depths_13),
    .io_inputs_depths_14(sltg_io_inputs_depths_14),
    .io_inputs_depths_15(sltg_io_inputs_depths_15),
    .io_inputs_depths_16(sltg_io_inputs_depths_16),
    .io_inputs_depths_17(sltg_io_inputs_depths_17),
    .io_inputs_depths_18(sltg_io_inputs_depths_18),
    .io_inputs_depths_19(sltg_io_inputs_depths_19),
    .io_inputs_depths_20(sltg_io_inputs_depths_20),
    .io_inputs_depths_21(sltg_io_inputs_depths_21),
    .io_inputs_depths_22(sltg_io_inputs_depths_22),
    .io_inputs_depths_23(sltg_io_inputs_depths_23),
    .io_inputs_depths_24(sltg_io_inputs_depths_24),
    .io_inputs_depths_25(sltg_io_inputs_depths_25),
    .io_inputs_depths_26(sltg_io_inputs_depths_26),
    .io_inputs_depths_27(sltg_io_inputs_depths_27),
    .io_inputs_depths_28(sltg_io_inputs_depths_28),
    .io_inputs_depths_29(sltg_io_inputs_depths_29),
    .io_inputs_depths_30(sltg_io_inputs_depths_30),
    .io_inputs_depths_31(sltg_io_inputs_depths_31),
    .io_inputs_validCharacters(sltg_io_inputs_validCharacters),
    .io_outputs_outputData_0(sltg_io_outputs_outputData_0),
    .io_outputs_outputData_1(sltg_io_outputs_outputData_1),
    .io_outputs_outputData_2(sltg_io_outputs_outputData_2),
    .io_outputs_outputData_3(sltg_io_outputs_outputData_3),
    .io_outputs_outputData_4(sltg_io_outputs_outputData_4),
    .io_outputs_outputData_5(sltg_io_outputs_outputData_5),
    .io_outputs_outputData_6(sltg_io_outputs_outputData_6),
    .io_outputs_outputData_7(sltg_io_outputs_outputData_7),
    .io_outputs_outputData_8(sltg_io_outputs_outputData_8),
    .io_outputs_outputData_9(sltg_io_outputs_outputData_9),
    .io_outputs_outputData_10(sltg_io_outputs_outputData_10),
    .io_outputs_outputData_11(sltg_io_outputs_outputData_11),
    .io_outputs_outputData_12(sltg_io_outputs_outputData_12),
    .io_outputs_outputData_13(sltg_io_outputs_outputData_13),
    .io_outputs_outputData_14(sltg_io_outputs_outputData_14),
    .io_outputs_outputData_15(sltg_io_outputs_outputData_15),
    .io_outputs_outputData_16(sltg_io_outputs_outputData_16),
    .io_outputs_outputData_17(sltg_io_outputs_outputData_17),
    .io_outputs_outputData_18(sltg_io_outputs_outputData_18),
    .io_outputs_outputData_19(sltg_io_outputs_outputData_19),
    .io_outputs_outputData_20(sltg_io_outputs_outputData_20),
    .io_outputs_outputData_21(sltg_io_outputs_outputData_21),
    .io_outputs_outputData_22(sltg_io_outputs_outputData_22),
    .io_outputs_outputData_23(sltg_io_outputs_outputData_23),
    .io_outputs_outputData_24(sltg_io_outputs_outputData_24),
    .io_outputs_outputData_25(sltg_io_outputs_outputData_25),
    .io_outputs_outputData_26(sltg_io_outputs_outputData_26),
    .io_outputs_outputData_27(sltg_io_outputs_outputData_27),
    .io_outputs_outputData_28(sltg_io_outputs_outputData_28),
    .io_outputs_outputData_29(sltg_io_outputs_outputData_29),
    .io_outputs_outputData_30(sltg_io_outputs_outputData_30),
    .io_outputs_outputData_31(sltg_io_outputs_outputData_31),
    .io_outputs_outputTags_0(sltg_io_outputs_outputTags_0),
    .io_outputs_outputTags_1(sltg_io_outputs_outputTags_1),
    .io_outputs_outputTags_2(sltg_io_outputs_outputTags_2),
    .io_outputs_outputTags_3(sltg_io_outputs_outputTags_3),
    .io_outputs_outputTags_4(sltg_io_outputs_outputTags_4),
    .io_outputs_outputTags_5(sltg_io_outputs_outputTags_5),
    .io_outputs_outputTags_6(sltg_io_outputs_outputTags_6),
    .io_outputs_outputTags_7(sltg_io_outputs_outputTags_7),
    .io_outputs_outputTags_8(sltg_io_outputs_outputTags_8),
    .io_outputs_outputTags_9(sltg_io_outputs_outputTags_9),
    .io_outputs_outputTags_10(sltg_io_outputs_outputTags_10),
    .io_outputs_outputTags_11(sltg_io_outputs_outputTags_11),
    .io_outputs_outputTags_12(sltg_io_outputs_outputTags_12),
    .io_outputs_outputTags_13(sltg_io_outputs_outputTags_13),
    .io_outputs_outputTags_14(sltg_io_outputs_outputTags_14),
    .io_outputs_outputTags_15(sltg_io_outputs_outputTags_15),
    .io_outputs_outputTags_16(sltg_io_outputs_outputTags_16),
    .io_outputs_outputTags_17(sltg_io_outputs_outputTags_17),
    .io_outputs_outputTags_18(sltg_io_outputs_outputTags_18),
    .io_outputs_outputTags_19(sltg_io_outputs_outputTags_19),
    .io_outputs_outputTags_20(sltg_io_outputs_outputTags_20),
    .io_outputs_outputTags_21(sltg_io_outputs_outputTags_21),
    .io_outputs_outputTags_22(sltg_io_outputs_outputTags_22),
    .io_outputs_outputTags_23(sltg_io_outputs_outputTags_23),
    .io_outputs_outputTags_24(sltg_io_outputs_outputTags_24),
    .io_outputs_outputTags_25(sltg_io_outputs_outputTags_25),
    .io_outputs_outputTags_26(sltg_io_outputs_outputTags_26),
    .io_outputs_outputTags_27(sltg_io_outputs_outputTags_27),
    .io_outputs_outputTags_28(sltg_io_outputs_outputTags_28),
    .io_outputs_outputTags_29(sltg_io_outputs_outputTags_29),
    .io_outputs_outputTags_30(sltg_io_outputs_outputTags_30),
    .io_outputs_outputTags_31(sltg_io_outputs_outputTags_31),
    .io_outputs_itemNumber(sltg_io_outputs_itemNumber),
    .io_finished(sltg_io_finished)
  );
  treeNormalizer tn ( // @[topLevel.scala 59:18]
    .clock(tn_clock),
    .reset(tn_reset),
    .io_start(tn_io_start),
    .io_inputs_outputData_0(tn_io_inputs_outputData_0),
    .io_inputs_outputData_1(tn_io_inputs_outputData_1),
    .io_inputs_outputData_2(tn_io_inputs_outputData_2),
    .io_inputs_outputData_3(tn_io_inputs_outputData_3),
    .io_inputs_outputData_4(tn_io_inputs_outputData_4),
    .io_inputs_outputData_5(tn_io_inputs_outputData_5),
    .io_inputs_outputData_6(tn_io_inputs_outputData_6),
    .io_inputs_outputData_7(tn_io_inputs_outputData_7),
    .io_inputs_outputData_8(tn_io_inputs_outputData_8),
    .io_inputs_outputData_9(tn_io_inputs_outputData_9),
    .io_inputs_outputData_10(tn_io_inputs_outputData_10),
    .io_inputs_outputData_11(tn_io_inputs_outputData_11),
    .io_inputs_outputData_12(tn_io_inputs_outputData_12),
    .io_inputs_outputData_13(tn_io_inputs_outputData_13),
    .io_inputs_outputData_14(tn_io_inputs_outputData_14),
    .io_inputs_outputData_15(tn_io_inputs_outputData_15),
    .io_inputs_outputData_16(tn_io_inputs_outputData_16),
    .io_inputs_outputData_17(tn_io_inputs_outputData_17),
    .io_inputs_outputData_18(tn_io_inputs_outputData_18),
    .io_inputs_outputData_19(tn_io_inputs_outputData_19),
    .io_inputs_outputData_20(tn_io_inputs_outputData_20),
    .io_inputs_outputData_21(tn_io_inputs_outputData_21),
    .io_inputs_outputData_22(tn_io_inputs_outputData_22),
    .io_inputs_outputData_23(tn_io_inputs_outputData_23),
    .io_inputs_outputData_24(tn_io_inputs_outputData_24),
    .io_inputs_outputData_25(tn_io_inputs_outputData_25),
    .io_inputs_outputData_26(tn_io_inputs_outputData_26),
    .io_inputs_outputData_27(tn_io_inputs_outputData_27),
    .io_inputs_outputData_28(tn_io_inputs_outputData_28),
    .io_inputs_outputData_29(tn_io_inputs_outputData_29),
    .io_inputs_outputData_30(tn_io_inputs_outputData_30),
    .io_inputs_outputData_31(tn_io_inputs_outputData_31),
    .io_inputs_outputTags_0(tn_io_inputs_outputTags_0),
    .io_inputs_outputTags_1(tn_io_inputs_outputTags_1),
    .io_inputs_outputTags_2(tn_io_inputs_outputTags_2),
    .io_inputs_outputTags_3(tn_io_inputs_outputTags_3),
    .io_inputs_outputTags_4(tn_io_inputs_outputTags_4),
    .io_inputs_outputTags_5(tn_io_inputs_outputTags_5),
    .io_inputs_outputTags_6(tn_io_inputs_outputTags_6),
    .io_inputs_outputTags_7(tn_io_inputs_outputTags_7),
    .io_inputs_outputTags_8(tn_io_inputs_outputTags_8),
    .io_inputs_outputTags_9(tn_io_inputs_outputTags_9),
    .io_inputs_outputTags_10(tn_io_inputs_outputTags_10),
    .io_inputs_outputTags_11(tn_io_inputs_outputTags_11),
    .io_inputs_outputTags_12(tn_io_inputs_outputTags_12),
    .io_inputs_outputTags_13(tn_io_inputs_outputTags_13),
    .io_inputs_outputTags_14(tn_io_inputs_outputTags_14),
    .io_inputs_outputTags_15(tn_io_inputs_outputTags_15),
    .io_inputs_outputTags_16(tn_io_inputs_outputTags_16),
    .io_inputs_outputTags_17(tn_io_inputs_outputTags_17),
    .io_inputs_outputTags_18(tn_io_inputs_outputTags_18),
    .io_inputs_outputTags_19(tn_io_inputs_outputTags_19),
    .io_inputs_outputTags_20(tn_io_inputs_outputTags_20),
    .io_inputs_outputTags_21(tn_io_inputs_outputTags_21),
    .io_inputs_outputTags_22(tn_io_inputs_outputTags_22),
    .io_inputs_outputTags_23(tn_io_inputs_outputTags_23),
    .io_inputs_outputTags_24(tn_io_inputs_outputTags_24),
    .io_inputs_outputTags_25(tn_io_inputs_outputTags_25),
    .io_inputs_outputTags_26(tn_io_inputs_outputTags_26),
    .io_inputs_outputTags_27(tn_io_inputs_outputTags_27),
    .io_inputs_outputTags_28(tn_io_inputs_outputTags_28),
    .io_inputs_outputTags_29(tn_io_inputs_outputTags_29),
    .io_inputs_outputTags_30(tn_io_inputs_outputTags_30),
    .io_inputs_outputTags_31(tn_io_inputs_outputTags_31),
    .io_inputs_itemNumber(tn_io_inputs_itemNumber),
    .io_outputs_charactersOut_0(tn_io_outputs_charactersOut_0),
    .io_outputs_charactersOut_1(tn_io_outputs_charactersOut_1),
    .io_outputs_charactersOut_2(tn_io_outputs_charactersOut_2),
    .io_outputs_charactersOut_3(tn_io_outputs_charactersOut_3),
    .io_outputs_charactersOut_4(tn_io_outputs_charactersOut_4),
    .io_outputs_charactersOut_5(tn_io_outputs_charactersOut_5),
    .io_outputs_charactersOut_6(tn_io_outputs_charactersOut_6),
    .io_outputs_charactersOut_7(tn_io_outputs_charactersOut_7),
    .io_outputs_charactersOut_8(tn_io_outputs_charactersOut_8),
    .io_outputs_charactersOut_9(tn_io_outputs_charactersOut_9),
    .io_outputs_charactersOut_10(tn_io_outputs_charactersOut_10),
    .io_outputs_charactersOut_11(tn_io_outputs_charactersOut_11),
    .io_outputs_charactersOut_12(tn_io_outputs_charactersOut_12),
    .io_outputs_charactersOut_13(tn_io_outputs_charactersOut_13),
    .io_outputs_charactersOut_14(tn_io_outputs_charactersOut_14),
    .io_outputs_charactersOut_15(tn_io_outputs_charactersOut_15),
    .io_outputs_charactersOut_16(tn_io_outputs_charactersOut_16),
    .io_outputs_charactersOut_17(tn_io_outputs_charactersOut_17),
    .io_outputs_charactersOut_18(tn_io_outputs_charactersOut_18),
    .io_outputs_charactersOut_19(tn_io_outputs_charactersOut_19),
    .io_outputs_charactersOut_20(tn_io_outputs_charactersOut_20),
    .io_outputs_charactersOut_21(tn_io_outputs_charactersOut_21),
    .io_outputs_charactersOut_22(tn_io_outputs_charactersOut_22),
    .io_outputs_charactersOut_23(tn_io_outputs_charactersOut_23),
    .io_outputs_charactersOut_24(tn_io_outputs_charactersOut_24),
    .io_outputs_charactersOut_25(tn_io_outputs_charactersOut_25),
    .io_outputs_charactersOut_26(tn_io_outputs_charactersOut_26),
    .io_outputs_charactersOut_27(tn_io_outputs_charactersOut_27),
    .io_outputs_charactersOut_28(tn_io_outputs_charactersOut_28),
    .io_outputs_charactersOut_29(tn_io_outputs_charactersOut_29),
    .io_outputs_charactersOut_30(tn_io_outputs_charactersOut_30),
    .io_outputs_charactersOut_31(tn_io_outputs_charactersOut_31),
    .io_outputs_depthsOut_0(tn_io_outputs_depthsOut_0),
    .io_outputs_depthsOut_1(tn_io_outputs_depthsOut_1),
    .io_outputs_depthsOut_2(tn_io_outputs_depthsOut_2),
    .io_outputs_depthsOut_3(tn_io_outputs_depthsOut_3),
    .io_outputs_depthsOut_4(tn_io_outputs_depthsOut_4),
    .io_outputs_depthsOut_5(tn_io_outputs_depthsOut_5),
    .io_outputs_depthsOut_6(tn_io_outputs_depthsOut_6),
    .io_outputs_depthsOut_7(tn_io_outputs_depthsOut_7),
    .io_outputs_depthsOut_8(tn_io_outputs_depthsOut_8),
    .io_outputs_depthsOut_9(tn_io_outputs_depthsOut_9),
    .io_outputs_depthsOut_10(tn_io_outputs_depthsOut_10),
    .io_outputs_depthsOut_11(tn_io_outputs_depthsOut_11),
    .io_outputs_depthsOut_12(tn_io_outputs_depthsOut_12),
    .io_outputs_depthsOut_13(tn_io_outputs_depthsOut_13),
    .io_outputs_depthsOut_14(tn_io_outputs_depthsOut_14),
    .io_outputs_depthsOut_15(tn_io_outputs_depthsOut_15),
    .io_outputs_depthsOut_16(tn_io_outputs_depthsOut_16),
    .io_outputs_depthsOut_17(tn_io_outputs_depthsOut_17),
    .io_outputs_depthsOut_18(tn_io_outputs_depthsOut_18),
    .io_outputs_depthsOut_19(tn_io_outputs_depthsOut_19),
    .io_outputs_depthsOut_20(tn_io_outputs_depthsOut_20),
    .io_outputs_depthsOut_21(tn_io_outputs_depthsOut_21),
    .io_outputs_depthsOut_22(tn_io_outputs_depthsOut_22),
    .io_outputs_depthsOut_23(tn_io_outputs_depthsOut_23),
    .io_outputs_depthsOut_24(tn_io_outputs_depthsOut_24),
    .io_outputs_depthsOut_25(tn_io_outputs_depthsOut_25),
    .io_outputs_depthsOut_26(tn_io_outputs_depthsOut_26),
    .io_outputs_depthsOut_27(tn_io_outputs_depthsOut_27),
    .io_outputs_depthsOut_28(tn_io_outputs_depthsOut_28),
    .io_outputs_depthsOut_29(tn_io_outputs_depthsOut_29),
    .io_outputs_depthsOut_30(tn_io_outputs_depthsOut_30),
    .io_outputs_depthsOut_31(tn_io_outputs_depthsOut_31),
    .io_outputs_validNodesOut(tn_io_outputs_validNodesOut),
    .io_finished(tn_io_finished)
  );
  codewordGenerator cg ( // @[topLevel.scala 69:18]
    .clock(cg_clock),
    .reset(cg_reset),
    .io_start(cg_io_start),
    .io_inputs_charactersOut_0(cg_io_inputs_charactersOut_0),
    .io_inputs_charactersOut_1(cg_io_inputs_charactersOut_1),
    .io_inputs_charactersOut_2(cg_io_inputs_charactersOut_2),
    .io_inputs_charactersOut_3(cg_io_inputs_charactersOut_3),
    .io_inputs_charactersOut_4(cg_io_inputs_charactersOut_4),
    .io_inputs_charactersOut_5(cg_io_inputs_charactersOut_5),
    .io_inputs_charactersOut_6(cg_io_inputs_charactersOut_6),
    .io_inputs_charactersOut_7(cg_io_inputs_charactersOut_7),
    .io_inputs_charactersOut_8(cg_io_inputs_charactersOut_8),
    .io_inputs_charactersOut_9(cg_io_inputs_charactersOut_9),
    .io_inputs_charactersOut_10(cg_io_inputs_charactersOut_10),
    .io_inputs_charactersOut_11(cg_io_inputs_charactersOut_11),
    .io_inputs_charactersOut_12(cg_io_inputs_charactersOut_12),
    .io_inputs_charactersOut_13(cg_io_inputs_charactersOut_13),
    .io_inputs_charactersOut_14(cg_io_inputs_charactersOut_14),
    .io_inputs_charactersOut_15(cg_io_inputs_charactersOut_15),
    .io_inputs_charactersOut_16(cg_io_inputs_charactersOut_16),
    .io_inputs_charactersOut_17(cg_io_inputs_charactersOut_17),
    .io_inputs_charactersOut_18(cg_io_inputs_charactersOut_18),
    .io_inputs_charactersOut_19(cg_io_inputs_charactersOut_19),
    .io_inputs_charactersOut_20(cg_io_inputs_charactersOut_20),
    .io_inputs_charactersOut_21(cg_io_inputs_charactersOut_21),
    .io_inputs_charactersOut_22(cg_io_inputs_charactersOut_22),
    .io_inputs_charactersOut_23(cg_io_inputs_charactersOut_23),
    .io_inputs_charactersOut_24(cg_io_inputs_charactersOut_24),
    .io_inputs_charactersOut_25(cg_io_inputs_charactersOut_25),
    .io_inputs_charactersOut_26(cg_io_inputs_charactersOut_26),
    .io_inputs_charactersOut_27(cg_io_inputs_charactersOut_27),
    .io_inputs_charactersOut_28(cg_io_inputs_charactersOut_28),
    .io_inputs_charactersOut_29(cg_io_inputs_charactersOut_29),
    .io_inputs_charactersOut_30(cg_io_inputs_charactersOut_30),
    .io_inputs_charactersOut_31(cg_io_inputs_charactersOut_31),
    .io_inputs_depthsOut_0(cg_io_inputs_depthsOut_0),
    .io_inputs_depthsOut_1(cg_io_inputs_depthsOut_1),
    .io_inputs_depthsOut_2(cg_io_inputs_depthsOut_2),
    .io_inputs_depthsOut_3(cg_io_inputs_depthsOut_3),
    .io_inputs_depthsOut_4(cg_io_inputs_depthsOut_4),
    .io_inputs_depthsOut_5(cg_io_inputs_depthsOut_5),
    .io_inputs_depthsOut_6(cg_io_inputs_depthsOut_6),
    .io_inputs_depthsOut_7(cg_io_inputs_depthsOut_7),
    .io_inputs_depthsOut_8(cg_io_inputs_depthsOut_8),
    .io_inputs_depthsOut_9(cg_io_inputs_depthsOut_9),
    .io_inputs_depthsOut_10(cg_io_inputs_depthsOut_10),
    .io_inputs_depthsOut_11(cg_io_inputs_depthsOut_11),
    .io_inputs_depthsOut_12(cg_io_inputs_depthsOut_12),
    .io_inputs_depthsOut_13(cg_io_inputs_depthsOut_13),
    .io_inputs_depthsOut_14(cg_io_inputs_depthsOut_14),
    .io_inputs_depthsOut_15(cg_io_inputs_depthsOut_15),
    .io_inputs_depthsOut_16(cg_io_inputs_depthsOut_16),
    .io_inputs_depthsOut_17(cg_io_inputs_depthsOut_17),
    .io_inputs_depthsOut_18(cg_io_inputs_depthsOut_18),
    .io_inputs_depthsOut_19(cg_io_inputs_depthsOut_19),
    .io_inputs_depthsOut_20(cg_io_inputs_depthsOut_20),
    .io_inputs_depthsOut_21(cg_io_inputs_depthsOut_21),
    .io_inputs_depthsOut_22(cg_io_inputs_depthsOut_22),
    .io_inputs_depthsOut_23(cg_io_inputs_depthsOut_23),
    .io_inputs_depthsOut_24(cg_io_inputs_depthsOut_24),
    .io_inputs_depthsOut_25(cg_io_inputs_depthsOut_25),
    .io_inputs_depthsOut_26(cg_io_inputs_depthsOut_26),
    .io_inputs_depthsOut_27(cg_io_inputs_depthsOut_27),
    .io_inputs_depthsOut_28(cg_io_inputs_depthsOut_28),
    .io_inputs_depthsOut_29(cg_io_inputs_depthsOut_29),
    .io_inputs_depthsOut_30(cg_io_inputs_depthsOut_30),
    .io_inputs_depthsOut_31(cg_io_inputs_depthsOut_31),
    .io_inputs_validNodesOut(cg_io_inputs_validNodesOut),
    .io_outputs_codewords_0(cg_io_outputs_codewords_0),
    .io_outputs_codewords_1(cg_io_outputs_codewords_1),
    .io_outputs_codewords_2(cg_io_outputs_codewords_2),
    .io_outputs_codewords_3(cg_io_outputs_codewords_3),
    .io_outputs_codewords_4(cg_io_outputs_codewords_4),
    .io_outputs_codewords_5(cg_io_outputs_codewords_5),
    .io_outputs_codewords_6(cg_io_outputs_codewords_6),
    .io_outputs_codewords_7(cg_io_outputs_codewords_7),
    .io_outputs_codewords_8(cg_io_outputs_codewords_8),
    .io_outputs_codewords_9(cg_io_outputs_codewords_9),
    .io_outputs_codewords_10(cg_io_outputs_codewords_10),
    .io_outputs_codewords_11(cg_io_outputs_codewords_11),
    .io_outputs_codewords_12(cg_io_outputs_codewords_12),
    .io_outputs_codewords_13(cg_io_outputs_codewords_13),
    .io_outputs_codewords_14(cg_io_outputs_codewords_14),
    .io_outputs_codewords_15(cg_io_outputs_codewords_15),
    .io_outputs_codewords_16(cg_io_outputs_codewords_16),
    .io_outputs_codewords_17(cg_io_outputs_codewords_17),
    .io_outputs_codewords_18(cg_io_outputs_codewords_18),
    .io_outputs_codewords_19(cg_io_outputs_codewords_19),
    .io_outputs_codewords_20(cg_io_outputs_codewords_20),
    .io_outputs_codewords_21(cg_io_outputs_codewords_21),
    .io_outputs_codewords_22(cg_io_outputs_codewords_22),
    .io_outputs_codewords_23(cg_io_outputs_codewords_23),
    .io_outputs_codewords_24(cg_io_outputs_codewords_24),
    .io_outputs_codewords_25(cg_io_outputs_codewords_25),
    .io_outputs_codewords_26(cg_io_outputs_codewords_26),
    .io_outputs_codewords_27(cg_io_outputs_codewords_27),
    .io_outputs_codewords_28(cg_io_outputs_codewords_28),
    .io_outputs_codewords_29(cg_io_outputs_codewords_29),
    .io_outputs_codewords_30(cg_io_outputs_codewords_30),
    .io_outputs_codewords_31(cg_io_outputs_codewords_31),
    .io_outputs_codewords_32(cg_io_outputs_codewords_32),
    .io_outputs_codewords_33(cg_io_outputs_codewords_33),
    .io_outputs_codewords_34(cg_io_outputs_codewords_34),
    .io_outputs_codewords_35(cg_io_outputs_codewords_35),
    .io_outputs_codewords_36(cg_io_outputs_codewords_36),
    .io_outputs_codewords_37(cg_io_outputs_codewords_37),
    .io_outputs_codewords_38(cg_io_outputs_codewords_38),
    .io_outputs_codewords_39(cg_io_outputs_codewords_39),
    .io_outputs_codewords_40(cg_io_outputs_codewords_40),
    .io_outputs_codewords_41(cg_io_outputs_codewords_41),
    .io_outputs_codewords_42(cg_io_outputs_codewords_42),
    .io_outputs_codewords_43(cg_io_outputs_codewords_43),
    .io_outputs_codewords_44(cg_io_outputs_codewords_44),
    .io_outputs_codewords_45(cg_io_outputs_codewords_45),
    .io_outputs_codewords_46(cg_io_outputs_codewords_46),
    .io_outputs_codewords_47(cg_io_outputs_codewords_47),
    .io_outputs_codewords_48(cg_io_outputs_codewords_48),
    .io_outputs_codewords_49(cg_io_outputs_codewords_49),
    .io_outputs_codewords_50(cg_io_outputs_codewords_50),
    .io_outputs_codewords_51(cg_io_outputs_codewords_51),
    .io_outputs_codewords_52(cg_io_outputs_codewords_52),
    .io_outputs_codewords_53(cg_io_outputs_codewords_53),
    .io_outputs_codewords_54(cg_io_outputs_codewords_54),
    .io_outputs_codewords_55(cg_io_outputs_codewords_55),
    .io_outputs_codewords_56(cg_io_outputs_codewords_56),
    .io_outputs_codewords_57(cg_io_outputs_codewords_57),
    .io_outputs_codewords_58(cg_io_outputs_codewords_58),
    .io_outputs_codewords_59(cg_io_outputs_codewords_59),
    .io_outputs_codewords_60(cg_io_outputs_codewords_60),
    .io_outputs_codewords_61(cg_io_outputs_codewords_61),
    .io_outputs_codewords_62(cg_io_outputs_codewords_62),
    .io_outputs_codewords_63(cg_io_outputs_codewords_63),
    .io_outputs_codewords_64(cg_io_outputs_codewords_64),
    .io_outputs_codewords_65(cg_io_outputs_codewords_65),
    .io_outputs_codewords_66(cg_io_outputs_codewords_66),
    .io_outputs_codewords_67(cg_io_outputs_codewords_67),
    .io_outputs_codewords_68(cg_io_outputs_codewords_68),
    .io_outputs_codewords_69(cg_io_outputs_codewords_69),
    .io_outputs_codewords_70(cg_io_outputs_codewords_70),
    .io_outputs_codewords_71(cg_io_outputs_codewords_71),
    .io_outputs_codewords_72(cg_io_outputs_codewords_72),
    .io_outputs_codewords_73(cg_io_outputs_codewords_73),
    .io_outputs_codewords_74(cg_io_outputs_codewords_74),
    .io_outputs_codewords_75(cg_io_outputs_codewords_75),
    .io_outputs_codewords_76(cg_io_outputs_codewords_76),
    .io_outputs_codewords_77(cg_io_outputs_codewords_77),
    .io_outputs_codewords_78(cg_io_outputs_codewords_78),
    .io_outputs_codewords_79(cg_io_outputs_codewords_79),
    .io_outputs_codewords_80(cg_io_outputs_codewords_80),
    .io_outputs_codewords_81(cg_io_outputs_codewords_81),
    .io_outputs_codewords_82(cg_io_outputs_codewords_82),
    .io_outputs_codewords_83(cg_io_outputs_codewords_83),
    .io_outputs_codewords_84(cg_io_outputs_codewords_84),
    .io_outputs_codewords_85(cg_io_outputs_codewords_85),
    .io_outputs_codewords_86(cg_io_outputs_codewords_86),
    .io_outputs_codewords_87(cg_io_outputs_codewords_87),
    .io_outputs_codewords_88(cg_io_outputs_codewords_88),
    .io_outputs_codewords_89(cg_io_outputs_codewords_89),
    .io_outputs_codewords_90(cg_io_outputs_codewords_90),
    .io_outputs_codewords_91(cg_io_outputs_codewords_91),
    .io_outputs_codewords_92(cg_io_outputs_codewords_92),
    .io_outputs_codewords_93(cg_io_outputs_codewords_93),
    .io_outputs_codewords_94(cg_io_outputs_codewords_94),
    .io_outputs_codewords_95(cg_io_outputs_codewords_95),
    .io_outputs_codewords_96(cg_io_outputs_codewords_96),
    .io_outputs_codewords_97(cg_io_outputs_codewords_97),
    .io_outputs_codewords_98(cg_io_outputs_codewords_98),
    .io_outputs_codewords_99(cg_io_outputs_codewords_99),
    .io_outputs_codewords_100(cg_io_outputs_codewords_100),
    .io_outputs_codewords_101(cg_io_outputs_codewords_101),
    .io_outputs_codewords_102(cg_io_outputs_codewords_102),
    .io_outputs_codewords_103(cg_io_outputs_codewords_103),
    .io_outputs_codewords_104(cg_io_outputs_codewords_104),
    .io_outputs_codewords_105(cg_io_outputs_codewords_105),
    .io_outputs_codewords_106(cg_io_outputs_codewords_106),
    .io_outputs_codewords_107(cg_io_outputs_codewords_107),
    .io_outputs_codewords_108(cg_io_outputs_codewords_108),
    .io_outputs_codewords_109(cg_io_outputs_codewords_109),
    .io_outputs_codewords_110(cg_io_outputs_codewords_110),
    .io_outputs_codewords_111(cg_io_outputs_codewords_111),
    .io_outputs_codewords_112(cg_io_outputs_codewords_112),
    .io_outputs_codewords_113(cg_io_outputs_codewords_113),
    .io_outputs_codewords_114(cg_io_outputs_codewords_114),
    .io_outputs_codewords_115(cg_io_outputs_codewords_115),
    .io_outputs_codewords_116(cg_io_outputs_codewords_116),
    .io_outputs_codewords_117(cg_io_outputs_codewords_117),
    .io_outputs_codewords_118(cg_io_outputs_codewords_118),
    .io_outputs_codewords_119(cg_io_outputs_codewords_119),
    .io_outputs_codewords_120(cg_io_outputs_codewords_120),
    .io_outputs_codewords_121(cg_io_outputs_codewords_121),
    .io_outputs_codewords_122(cg_io_outputs_codewords_122),
    .io_outputs_codewords_123(cg_io_outputs_codewords_123),
    .io_outputs_codewords_124(cg_io_outputs_codewords_124),
    .io_outputs_codewords_125(cg_io_outputs_codewords_125),
    .io_outputs_codewords_126(cg_io_outputs_codewords_126),
    .io_outputs_codewords_127(cg_io_outputs_codewords_127),
    .io_outputs_codewords_128(cg_io_outputs_codewords_128),
    .io_outputs_codewords_129(cg_io_outputs_codewords_129),
    .io_outputs_codewords_130(cg_io_outputs_codewords_130),
    .io_outputs_codewords_131(cg_io_outputs_codewords_131),
    .io_outputs_codewords_132(cg_io_outputs_codewords_132),
    .io_outputs_codewords_133(cg_io_outputs_codewords_133),
    .io_outputs_codewords_134(cg_io_outputs_codewords_134),
    .io_outputs_codewords_135(cg_io_outputs_codewords_135),
    .io_outputs_codewords_136(cg_io_outputs_codewords_136),
    .io_outputs_codewords_137(cg_io_outputs_codewords_137),
    .io_outputs_codewords_138(cg_io_outputs_codewords_138),
    .io_outputs_codewords_139(cg_io_outputs_codewords_139),
    .io_outputs_codewords_140(cg_io_outputs_codewords_140),
    .io_outputs_codewords_141(cg_io_outputs_codewords_141),
    .io_outputs_codewords_142(cg_io_outputs_codewords_142),
    .io_outputs_codewords_143(cg_io_outputs_codewords_143),
    .io_outputs_codewords_144(cg_io_outputs_codewords_144),
    .io_outputs_codewords_145(cg_io_outputs_codewords_145),
    .io_outputs_codewords_146(cg_io_outputs_codewords_146),
    .io_outputs_codewords_147(cg_io_outputs_codewords_147),
    .io_outputs_codewords_148(cg_io_outputs_codewords_148),
    .io_outputs_codewords_149(cg_io_outputs_codewords_149),
    .io_outputs_codewords_150(cg_io_outputs_codewords_150),
    .io_outputs_codewords_151(cg_io_outputs_codewords_151),
    .io_outputs_codewords_152(cg_io_outputs_codewords_152),
    .io_outputs_codewords_153(cg_io_outputs_codewords_153),
    .io_outputs_codewords_154(cg_io_outputs_codewords_154),
    .io_outputs_codewords_155(cg_io_outputs_codewords_155),
    .io_outputs_codewords_156(cg_io_outputs_codewords_156),
    .io_outputs_codewords_157(cg_io_outputs_codewords_157),
    .io_outputs_codewords_158(cg_io_outputs_codewords_158),
    .io_outputs_codewords_159(cg_io_outputs_codewords_159),
    .io_outputs_codewords_160(cg_io_outputs_codewords_160),
    .io_outputs_codewords_161(cg_io_outputs_codewords_161),
    .io_outputs_codewords_162(cg_io_outputs_codewords_162),
    .io_outputs_codewords_163(cg_io_outputs_codewords_163),
    .io_outputs_codewords_164(cg_io_outputs_codewords_164),
    .io_outputs_codewords_165(cg_io_outputs_codewords_165),
    .io_outputs_codewords_166(cg_io_outputs_codewords_166),
    .io_outputs_codewords_167(cg_io_outputs_codewords_167),
    .io_outputs_codewords_168(cg_io_outputs_codewords_168),
    .io_outputs_codewords_169(cg_io_outputs_codewords_169),
    .io_outputs_codewords_170(cg_io_outputs_codewords_170),
    .io_outputs_codewords_171(cg_io_outputs_codewords_171),
    .io_outputs_codewords_172(cg_io_outputs_codewords_172),
    .io_outputs_codewords_173(cg_io_outputs_codewords_173),
    .io_outputs_codewords_174(cg_io_outputs_codewords_174),
    .io_outputs_codewords_175(cg_io_outputs_codewords_175),
    .io_outputs_codewords_176(cg_io_outputs_codewords_176),
    .io_outputs_codewords_177(cg_io_outputs_codewords_177),
    .io_outputs_codewords_178(cg_io_outputs_codewords_178),
    .io_outputs_codewords_179(cg_io_outputs_codewords_179),
    .io_outputs_codewords_180(cg_io_outputs_codewords_180),
    .io_outputs_codewords_181(cg_io_outputs_codewords_181),
    .io_outputs_codewords_182(cg_io_outputs_codewords_182),
    .io_outputs_codewords_183(cg_io_outputs_codewords_183),
    .io_outputs_codewords_184(cg_io_outputs_codewords_184),
    .io_outputs_codewords_185(cg_io_outputs_codewords_185),
    .io_outputs_codewords_186(cg_io_outputs_codewords_186),
    .io_outputs_codewords_187(cg_io_outputs_codewords_187),
    .io_outputs_codewords_188(cg_io_outputs_codewords_188),
    .io_outputs_codewords_189(cg_io_outputs_codewords_189),
    .io_outputs_codewords_190(cg_io_outputs_codewords_190),
    .io_outputs_codewords_191(cg_io_outputs_codewords_191),
    .io_outputs_codewords_192(cg_io_outputs_codewords_192),
    .io_outputs_codewords_193(cg_io_outputs_codewords_193),
    .io_outputs_codewords_194(cg_io_outputs_codewords_194),
    .io_outputs_codewords_195(cg_io_outputs_codewords_195),
    .io_outputs_codewords_196(cg_io_outputs_codewords_196),
    .io_outputs_codewords_197(cg_io_outputs_codewords_197),
    .io_outputs_codewords_198(cg_io_outputs_codewords_198),
    .io_outputs_codewords_199(cg_io_outputs_codewords_199),
    .io_outputs_codewords_200(cg_io_outputs_codewords_200),
    .io_outputs_codewords_201(cg_io_outputs_codewords_201),
    .io_outputs_codewords_202(cg_io_outputs_codewords_202),
    .io_outputs_codewords_203(cg_io_outputs_codewords_203),
    .io_outputs_codewords_204(cg_io_outputs_codewords_204),
    .io_outputs_codewords_205(cg_io_outputs_codewords_205),
    .io_outputs_codewords_206(cg_io_outputs_codewords_206),
    .io_outputs_codewords_207(cg_io_outputs_codewords_207),
    .io_outputs_codewords_208(cg_io_outputs_codewords_208),
    .io_outputs_codewords_209(cg_io_outputs_codewords_209),
    .io_outputs_codewords_210(cg_io_outputs_codewords_210),
    .io_outputs_codewords_211(cg_io_outputs_codewords_211),
    .io_outputs_codewords_212(cg_io_outputs_codewords_212),
    .io_outputs_codewords_213(cg_io_outputs_codewords_213),
    .io_outputs_codewords_214(cg_io_outputs_codewords_214),
    .io_outputs_codewords_215(cg_io_outputs_codewords_215),
    .io_outputs_codewords_216(cg_io_outputs_codewords_216),
    .io_outputs_codewords_217(cg_io_outputs_codewords_217),
    .io_outputs_codewords_218(cg_io_outputs_codewords_218),
    .io_outputs_codewords_219(cg_io_outputs_codewords_219),
    .io_outputs_codewords_220(cg_io_outputs_codewords_220),
    .io_outputs_codewords_221(cg_io_outputs_codewords_221),
    .io_outputs_codewords_222(cg_io_outputs_codewords_222),
    .io_outputs_codewords_223(cg_io_outputs_codewords_223),
    .io_outputs_codewords_224(cg_io_outputs_codewords_224),
    .io_outputs_codewords_225(cg_io_outputs_codewords_225),
    .io_outputs_codewords_226(cg_io_outputs_codewords_226),
    .io_outputs_codewords_227(cg_io_outputs_codewords_227),
    .io_outputs_codewords_228(cg_io_outputs_codewords_228),
    .io_outputs_codewords_229(cg_io_outputs_codewords_229),
    .io_outputs_codewords_230(cg_io_outputs_codewords_230),
    .io_outputs_codewords_231(cg_io_outputs_codewords_231),
    .io_outputs_codewords_232(cg_io_outputs_codewords_232),
    .io_outputs_codewords_233(cg_io_outputs_codewords_233),
    .io_outputs_codewords_234(cg_io_outputs_codewords_234),
    .io_outputs_codewords_235(cg_io_outputs_codewords_235),
    .io_outputs_codewords_236(cg_io_outputs_codewords_236),
    .io_outputs_codewords_237(cg_io_outputs_codewords_237),
    .io_outputs_codewords_238(cg_io_outputs_codewords_238),
    .io_outputs_codewords_239(cg_io_outputs_codewords_239),
    .io_outputs_codewords_240(cg_io_outputs_codewords_240),
    .io_outputs_codewords_241(cg_io_outputs_codewords_241),
    .io_outputs_codewords_242(cg_io_outputs_codewords_242),
    .io_outputs_codewords_243(cg_io_outputs_codewords_243),
    .io_outputs_codewords_244(cg_io_outputs_codewords_244),
    .io_outputs_codewords_245(cg_io_outputs_codewords_245),
    .io_outputs_codewords_246(cg_io_outputs_codewords_246),
    .io_outputs_codewords_247(cg_io_outputs_codewords_247),
    .io_outputs_codewords_248(cg_io_outputs_codewords_248),
    .io_outputs_codewords_249(cg_io_outputs_codewords_249),
    .io_outputs_codewords_250(cg_io_outputs_codewords_250),
    .io_outputs_codewords_251(cg_io_outputs_codewords_251),
    .io_outputs_codewords_252(cg_io_outputs_codewords_252),
    .io_outputs_codewords_253(cg_io_outputs_codewords_253),
    .io_outputs_codewords_254(cg_io_outputs_codewords_254),
    .io_outputs_codewords_255(cg_io_outputs_codewords_255),
    .io_outputs_lengths_0(cg_io_outputs_lengths_0),
    .io_outputs_lengths_1(cg_io_outputs_lengths_1),
    .io_outputs_lengths_2(cg_io_outputs_lengths_2),
    .io_outputs_lengths_3(cg_io_outputs_lengths_3),
    .io_outputs_lengths_4(cg_io_outputs_lengths_4),
    .io_outputs_lengths_5(cg_io_outputs_lengths_5),
    .io_outputs_lengths_6(cg_io_outputs_lengths_6),
    .io_outputs_lengths_7(cg_io_outputs_lengths_7),
    .io_outputs_lengths_8(cg_io_outputs_lengths_8),
    .io_outputs_lengths_9(cg_io_outputs_lengths_9),
    .io_outputs_lengths_10(cg_io_outputs_lengths_10),
    .io_outputs_lengths_11(cg_io_outputs_lengths_11),
    .io_outputs_lengths_12(cg_io_outputs_lengths_12),
    .io_outputs_lengths_13(cg_io_outputs_lengths_13),
    .io_outputs_lengths_14(cg_io_outputs_lengths_14),
    .io_outputs_lengths_15(cg_io_outputs_lengths_15),
    .io_outputs_lengths_16(cg_io_outputs_lengths_16),
    .io_outputs_lengths_17(cg_io_outputs_lengths_17),
    .io_outputs_lengths_18(cg_io_outputs_lengths_18),
    .io_outputs_lengths_19(cg_io_outputs_lengths_19),
    .io_outputs_lengths_20(cg_io_outputs_lengths_20),
    .io_outputs_lengths_21(cg_io_outputs_lengths_21),
    .io_outputs_lengths_22(cg_io_outputs_lengths_22),
    .io_outputs_lengths_23(cg_io_outputs_lengths_23),
    .io_outputs_lengths_24(cg_io_outputs_lengths_24),
    .io_outputs_lengths_25(cg_io_outputs_lengths_25),
    .io_outputs_lengths_26(cg_io_outputs_lengths_26),
    .io_outputs_lengths_27(cg_io_outputs_lengths_27),
    .io_outputs_lengths_28(cg_io_outputs_lengths_28),
    .io_outputs_lengths_29(cg_io_outputs_lengths_29),
    .io_outputs_lengths_30(cg_io_outputs_lengths_30),
    .io_outputs_lengths_31(cg_io_outputs_lengths_31),
    .io_outputs_lengths_32(cg_io_outputs_lengths_32),
    .io_outputs_lengths_33(cg_io_outputs_lengths_33),
    .io_outputs_lengths_34(cg_io_outputs_lengths_34),
    .io_outputs_lengths_35(cg_io_outputs_lengths_35),
    .io_outputs_lengths_36(cg_io_outputs_lengths_36),
    .io_outputs_lengths_37(cg_io_outputs_lengths_37),
    .io_outputs_lengths_38(cg_io_outputs_lengths_38),
    .io_outputs_lengths_39(cg_io_outputs_lengths_39),
    .io_outputs_lengths_40(cg_io_outputs_lengths_40),
    .io_outputs_lengths_41(cg_io_outputs_lengths_41),
    .io_outputs_lengths_42(cg_io_outputs_lengths_42),
    .io_outputs_lengths_43(cg_io_outputs_lengths_43),
    .io_outputs_lengths_44(cg_io_outputs_lengths_44),
    .io_outputs_lengths_45(cg_io_outputs_lengths_45),
    .io_outputs_lengths_46(cg_io_outputs_lengths_46),
    .io_outputs_lengths_47(cg_io_outputs_lengths_47),
    .io_outputs_lengths_48(cg_io_outputs_lengths_48),
    .io_outputs_lengths_49(cg_io_outputs_lengths_49),
    .io_outputs_lengths_50(cg_io_outputs_lengths_50),
    .io_outputs_lengths_51(cg_io_outputs_lengths_51),
    .io_outputs_lengths_52(cg_io_outputs_lengths_52),
    .io_outputs_lengths_53(cg_io_outputs_lengths_53),
    .io_outputs_lengths_54(cg_io_outputs_lengths_54),
    .io_outputs_lengths_55(cg_io_outputs_lengths_55),
    .io_outputs_lengths_56(cg_io_outputs_lengths_56),
    .io_outputs_lengths_57(cg_io_outputs_lengths_57),
    .io_outputs_lengths_58(cg_io_outputs_lengths_58),
    .io_outputs_lengths_59(cg_io_outputs_lengths_59),
    .io_outputs_lengths_60(cg_io_outputs_lengths_60),
    .io_outputs_lengths_61(cg_io_outputs_lengths_61),
    .io_outputs_lengths_62(cg_io_outputs_lengths_62),
    .io_outputs_lengths_63(cg_io_outputs_lengths_63),
    .io_outputs_lengths_64(cg_io_outputs_lengths_64),
    .io_outputs_lengths_65(cg_io_outputs_lengths_65),
    .io_outputs_lengths_66(cg_io_outputs_lengths_66),
    .io_outputs_lengths_67(cg_io_outputs_lengths_67),
    .io_outputs_lengths_68(cg_io_outputs_lengths_68),
    .io_outputs_lengths_69(cg_io_outputs_lengths_69),
    .io_outputs_lengths_70(cg_io_outputs_lengths_70),
    .io_outputs_lengths_71(cg_io_outputs_lengths_71),
    .io_outputs_lengths_72(cg_io_outputs_lengths_72),
    .io_outputs_lengths_73(cg_io_outputs_lengths_73),
    .io_outputs_lengths_74(cg_io_outputs_lengths_74),
    .io_outputs_lengths_75(cg_io_outputs_lengths_75),
    .io_outputs_lengths_76(cg_io_outputs_lengths_76),
    .io_outputs_lengths_77(cg_io_outputs_lengths_77),
    .io_outputs_lengths_78(cg_io_outputs_lengths_78),
    .io_outputs_lengths_79(cg_io_outputs_lengths_79),
    .io_outputs_lengths_80(cg_io_outputs_lengths_80),
    .io_outputs_lengths_81(cg_io_outputs_lengths_81),
    .io_outputs_lengths_82(cg_io_outputs_lengths_82),
    .io_outputs_lengths_83(cg_io_outputs_lengths_83),
    .io_outputs_lengths_84(cg_io_outputs_lengths_84),
    .io_outputs_lengths_85(cg_io_outputs_lengths_85),
    .io_outputs_lengths_86(cg_io_outputs_lengths_86),
    .io_outputs_lengths_87(cg_io_outputs_lengths_87),
    .io_outputs_lengths_88(cg_io_outputs_lengths_88),
    .io_outputs_lengths_89(cg_io_outputs_lengths_89),
    .io_outputs_lengths_90(cg_io_outputs_lengths_90),
    .io_outputs_lengths_91(cg_io_outputs_lengths_91),
    .io_outputs_lengths_92(cg_io_outputs_lengths_92),
    .io_outputs_lengths_93(cg_io_outputs_lengths_93),
    .io_outputs_lengths_94(cg_io_outputs_lengths_94),
    .io_outputs_lengths_95(cg_io_outputs_lengths_95),
    .io_outputs_lengths_96(cg_io_outputs_lengths_96),
    .io_outputs_lengths_97(cg_io_outputs_lengths_97),
    .io_outputs_lengths_98(cg_io_outputs_lengths_98),
    .io_outputs_lengths_99(cg_io_outputs_lengths_99),
    .io_outputs_lengths_100(cg_io_outputs_lengths_100),
    .io_outputs_lengths_101(cg_io_outputs_lengths_101),
    .io_outputs_lengths_102(cg_io_outputs_lengths_102),
    .io_outputs_lengths_103(cg_io_outputs_lengths_103),
    .io_outputs_lengths_104(cg_io_outputs_lengths_104),
    .io_outputs_lengths_105(cg_io_outputs_lengths_105),
    .io_outputs_lengths_106(cg_io_outputs_lengths_106),
    .io_outputs_lengths_107(cg_io_outputs_lengths_107),
    .io_outputs_lengths_108(cg_io_outputs_lengths_108),
    .io_outputs_lengths_109(cg_io_outputs_lengths_109),
    .io_outputs_lengths_110(cg_io_outputs_lengths_110),
    .io_outputs_lengths_111(cg_io_outputs_lengths_111),
    .io_outputs_lengths_112(cg_io_outputs_lengths_112),
    .io_outputs_lengths_113(cg_io_outputs_lengths_113),
    .io_outputs_lengths_114(cg_io_outputs_lengths_114),
    .io_outputs_lengths_115(cg_io_outputs_lengths_115),
    .io_outputs_lengths_116(cg_io_outputs_lengths_116),
    .io_outputs_lengths_117(cg_io_outputs_lengths_117),
    .io_outputs_lengths_118(cg_io_outputs_lengths_118),
    .io_outputs_lengths_119(cg_io_outputs_lengths_119),
    .io_outputs_lengths_120(cg_io_outputs_lengths_120),
    .io_outputs_lengths_121(cg_io_outputs_lengths_121),
    .io_outputs_lengths_122(cg_io_outputs_lengths_122),
    .io_outputs_lengths_123(cg_io_outputs_lengths_123),
    .io_outputs_lengths_124(cg_io_outputs_lengths_124),
    .io_outputs_lengths_125(cg_io_outputs_lengths_125),
    .io_outputs_lengths_126(cg_io_outputs_lengths_126),
    .io_outputs_lengths_127(cg_io_outputs_lengths_127),
    .io_outputs_lengths_128(cg_io_outputs_lengths_128),
    .io_outputs_lengths_129(cg_io_outputs_lengths_129),
    .io_outputs_lengths_130(cg_io_outputs_lengths_130),
    .io_outputs_lengths_131(cg_io_outputs_lengths_131),
    .io_outputs_lengths_132(cg_io_outputs_lengths_132),
    .io_outputs_lengths_133(cg_io_outputs_lengths_133),
    .io_outputs_lengths_134(cg_io_outputs_lengths_134),
    .io_outputs_lengths_135(cg_io_outputs_lengths_135),
    .io_outputs_lengths_136(cg_io_outputs_lengths_136),
    .io_outputs_lengths_137(cg_io_outputs_lengths_137),
    .io_outputs_lengths_138(cg_io_outputs_lengths_138),
    .io_outputs_lengths_139(cg_io_outputs_lengths_139),
    .io_outputs_lengths_140(cg_io_outputs_lengths_140),
    .io_outputs_lengths_141(cg_io_outputs_lengths_141),
    .io_outputs_lengths_142(cg_io_outputs_lengths_142),
    .io_outputs_lengths_143(cg_io_outputs_lengths_143),
    .io_outputs_lengths_144(cg_io_outputs_lengths_144),
    .io_outputs_lengths_145(cg_io_outputs_lengths_145),
    .io_outputs_lengths_146(cg_io_outputs_lengths_146),
    .io_outputs_lengths_147(cg_io_outputs_lengths_147),
    .io_outputs_lengths_148(cg_io_outputs_lengths_148),
    .io_outputs_lengths_149(cg_io_outputs_lengths_149),
    .io_outputs_lengths_150(cg_io_outputs_lengths_150),
    .io_outputs_lengths_151(cg_io_outputs_lengths_151),
    .io_outputs_lengths_152(cg_io_outputs_lengths_152),
    .io_outputs_lengths_153(cg_io_outputs_lengths_153),
    .io_outputs_lengths_154(cg_io_outputs_lengths_154),
    .io_outputs_lengths_155(cg_io_outputs_lengths_155),
    .io_outputs_lengths_156(cg_io_outputs_lengths_156),
    .io_outputs_lengths_157(cg_io_outputs_lengths_157),
    .io_outputs_lengths_158(cg_io_outputs_lengths_158),
    .io_outputs_lengths_159(cg_io_outputs_lengths_159),
    .io_outputs_lengths_160(cg_io_outputs_lengths_160),
    .io_outputs_lengths_161(cg_io_outputs_lengths_161),
    .io_outputs_lengths_162(cg_io_outputs_lengths_162),
    .io_outputs_lengths_163(cg_io_outputs_lengths_163),
    .io_outputs_lengths_164(cg_io_outputs_lengths_164),
    .io_outputs_lengths_165(cg_io_outputs_lengths_165),
    .io_outputs_lengths_166(cg_io_outputs_lengths_166),
    .io_outputs_lengths_167(cg_io_outputs_lengths_167),
    .io_outputs_lengths_168(cg_io_outputs_lengths_168),
    .io_outputs_lengths_169(cg_io_outputs_lengths_169),
    .io_outputs_lengths_170(cg_io_outputs_lengths_170),
    .io_outputs_lengths_171(cg_io_outputs_lengths_171),
    .io_outputs_lengths_172(cg_io_outputs_lengths_172),
    .io_outputs_lengths_173(cg_io_outputs_lengths_173),
    .io_outputs_lengths_174(cg_io_outputs_lengths_174),
    .io_outputs_lengths_175(cg_io_outputs_lengths_175),
    .io_outputs_lengths_176(cg_io_outputs_lengths_176),
    .io_outputs_lengths_177(cg_io_outputs_lengths_177),
    .io_outputs_lengths_178(cg_io_outputs_lengths_178),
    .io_outputs_lengths_179(cg_io_outputs_lengths_179),
    .io_outputs_lengths_180(cg_io_outputs_lengths_180),
    .io_outputs_lengths_181(cg_io_outputs_lengths_181),
    .io_outputs_lengths_182(cg_io_outputs_lengths_182),
    .io_outputs_lengths_183(cg_io_outputs_lengths_183),
    .io_outputs_lengths_184(cg_io_outputs_lengths_184),
    .io_outputs_lengths_185(cg_io_outputs_lengths_185),
    .io_outputs_lengths_186(cg_io_outputs_lengths_186),
    .io_outputs_lengths_187(cg_io_outputs_lengths_187),
    .io_outputs_lengths_188(cg_io_outputs_lengths_188),
    .io_outputs_lengths_189(cg_io_outputs_lengths_189),
    .io_outputs_lengths_190(cg_io_outputs_lengths_190),
    .io_outputs_lengths_191(cg_io_outputs_lengths_191),
    .io_outputs_lengths_192(cg_io_outputs_lengths_192),
    .io_outputs_lengths_193(cg_io_outputs_lengths_193),
    .io_outputs_lengths_194(cg_io_outputs_lengths_194),
    .io_outputs_lengths_195(cg_io_outputs_lengths_195),
    .io_outputs_lengths_196(cg_io_outputs_lengths_196),
    .io_outputs_lengths_197(cg_io_outputs_lengths_197),
    .io_outputs_lengths_198(cg_io_outputs_lengths_198),
    .io_outputs_lengths_199(cg_io_outputs_lengths_199),
    .io_outputs_lengths_200(cg_io_outputs_lengths_200),
    .io_outputs_lengths_201(cg_io_outputs_lengths_201),
    .io_outputs_lengths_202(cg_io_outputs_lengths_202),
    .io_outputs_lengths_203(cg_io_outputs_lengths_203),
    .io_outputs_lengths_204(cg_io_outputs_lengths_204),
    .io_outputs_lengths_205(cg_io_outputs_lengths_205),
    .io_outputs_lengths_206(cg_io_outputs_lengths_206),
    .io_outputs_lengths_207(cg_io_outputs_lengths_207),
    .io_outputs_lengths_208(cg_io_outputs_lengths_208),
    .io_outputs_lengths_209(cg_io_outputs_lengths_209),
    .io_outputs_lengths_210(cg_io_outputs_lengths_210),
    .io_outputs_lengths_211(cg_io_outputs_lengths_211),
    .io_outputs_lengths_212(cg_io_outputs_lengths_212),
    .io_outputs_lengths_213(cg_io_outputs_lengths_213),
    .io_outputs_lengths_214(cg_io_outputs_lengths_214),
    .io_outputs_lengths_215(cg_io_outputs_lengths_215),
    .io_outputs_lengths_216(cg_io_outputs_lengths_216),
    .io_outputs_lengths_217(cg_io_outputs_lengths_217),
    .io_outputs_lengths_218(cg_io_outputs_lengths_218),
    .io_outputs_lengths_219(cg_io_outputs_lengths_219),
    .io_outputs_lengths_220(cg_io_outputs_lengths_220),
    .io_outputs_lengths_221(cg_io_outputs_lengths_221),
    .io_outputs_lengths_222(cg_io_outputs_lengths_222),
    .io_outputs_lengths_223(cg_io_outputs_lengths_223),
    .io_outputs_lengths_224(cg_io_outputs_lengths_224),
    .io_outputs_lengths_225(cg_io_outputs_lengths_225),
    .io_outputs_lengths_226(cg_io_outputs_lengths_226),
    .io_outputs_lengths_227(cg_io_outputs_lengths_227),
    .io_outputs_lengths_228(cg_io_outputs_lengths_228),
    .io_outputs_lengths_229(cg_io_outputs_lengths_229),
    .io_outputs_lengths_230(cg_io_outputs_lengths_230),
    .io_outputs_lengths_231(cg_io_outputs_lengths_231),
    .io_outputs_lengths_232(cg_io_outputs_lengths_232),
    .io_outputs_lengths_233(cg_io_outputs_lengths_233),
    .io_outputs_lengths_234(cg_io_outputs_lengths_234),
    .io_outputs_lengths_235(cg_io_outputs_lengths_235),
    .io_outputs_lengths_236(cg_io_outputs_lengths_236),
    .io_outputs_lengths_237(cg_io_outputs_lengths_237),
    .io_outputs_lengths_238(cg_io_outputs_lengths_238),
    .io_outputs_lengths_239(cg_io_outputs_lengths_239),
    .io_outputs_lengths_240(cg_io_outputs_lengths_240),
    .io_outputs_lengths_241(cg_io_outputs_lengths_241),
    .io_outputs_lengths_242(cg_io_outputs_lengths_242),
    .io_outputs_lengths_243(cg_io_outputs_lengths_243),
    .io_outputs_lengths_244(cg_io_outputs_lengths_244),
    .io_outputs_lengths_245(cg_io_outputs_lengths_245),
    .io_outputs_lengths_246(cg_io_outputs_lengths_246),
    .io_outputs_lengths_247(cg_io_outputs_lengths_247),
    .io_outputs_lengths_248(cg_io_outputs_lengths_248),
    .io_outputs_lengths_249(cg_io_outputs_lengths_249),
    .io_outputs_lengths_250(cg_io_outputs_lengths_250),
    .io_outputs_lengths_251(cg_io_outputs_lengths_251),
    .io_outputs_lengths_252(cg_io_outputs_lengths_252),
    .io_outputs_lengths_253(cg_io_outputs_lengths_253),
    .io_outputs_lengths_254(cg_io_outputs_lengths_254),
    .io_outputs_lengths_255(cg_io_outputs_lengths_255),
    .io_outputs_charactersOut_0(cg_io_outputs_charactersOut_0),
    .io_outputs_charactersOut_1(cg_io_outputs_charactersOut_1),
    .io_outputs_charactersOut_2(cg_io_outputs_charactersOut_2),
    .io_outputs_charactersOut_3(cg_io_outputs_charactersOut_3),
    .io_outputs_charactersOut_4(cg_io_outputs_charactersOut_4),
    .io_outputs_charactersOut_5(cg_io_outputs_charactersOut_5),
    .io_outputs_charactersOut_6(cg_io_outputs_charactersOut_6),
    .io_outputs_charactersOut_7(cg_io_outputs_charactersOut_7),
    .io_outputs_charactersOut_8(cg_io_outputs_charactersOut_8),
    .io_outputs_charactersOut_9(cg_io_outputs_charactersOut_9),
    .io_outputs_charactersOut_10(cg_io_outputs_charactersOut_10),
    .io_outputs_charactersOut_11(cg_io_outputs_charactersOut_11),
    .io_outputs_charactersOut_12(cg_io_outputs_charactersOut_12),
    .io_outputs_charactersOut_13(cg_io_outputs_charactersOut_13),
    .io_outputs_charactersOut_14(cg_io_outputs_charactersOut_14),
    .io_outputs_charactersOut_15(cg_io_outputs_charactersOut_15),
    .io_outputs_charactersOut_16(cg_io_outputs_charactersOut_16),
    .io_outputs_charactersOut_17(cg_io_outputs_charactersOut_17),
    .io_outputs_charactersOut_18(cg_io_outputs_charactersOut_18),
    .io_outputs_charactersOut_19(cg_io_outputs_charactersOut_19),
    .io_outputs_charactersOut_20(cg_io_outputs_charactersOut_20),
    .io_outputs_charactersOut_21(cg_io_outputs_charactersOut_21),
    .io_outputs_charactersOut_22(cg_io_outputs_charactersOut_22),
    .io_outputs_charactersOut_23(cg_io_outputs_charactersOut_23),
    .io_outputs_charactersOut_24(cg_io_outputs_charactersOut_24),
    .io_outputs_charactersOut_25(cg_io_outputs_charactersOut_25),
    .io_outputs_charactersOut_26(cg_io_outputs_charactersOut_26),
    .io_outputs_charactersOut_27(cg_io_outputs_charactersOut_27),
    .io_outputs_charactersOut_28(cg_io_outputs_charactersOut_28),
    .io_outputs_charactersOut_29(cg_io_outputs_charactersOut_29),
    .io_outputs_charactersOut_30(cg_io_outputs_charactersOut_30),
    .io_outputs_charactersOut_31(cg_io_outputs_charactersOut_31),
    .io_outputs_nodes(cg_io_outputs_nodes),
    .io_outputs_escapeCharacterLength(cg_io_outputs_escapeCharacterLength),
    .io_outputs_escapeCodeword(cg_io_outputs_escapeCodeword),
    .io_finished(cg_io_finished)
  );
  compressorOutput co ( // @[topLevel.scala 72:18]
    .clock(co_clock),
    .reset(co_reset),
    .io_start(co_io_start),
    .io_dataIn_0_currentByteOut(co_io_dataIn_0_currentByteOut),
    .io_dataIn_0_dataIn_0(co_io_dataIn_0_dataIn_0),
    .io_dataIn_0_valid(co_io_dataIn_0_valid),
    .io_dataIn_0_ready(co_io_dataIn_0_ready),
    .io_inputs_codewords_0(co_io_inputs_codewords_0),
    .io_inputs_codewords_1(co_io_inputs_codewords_1),
    .io_inputs_codewords_2(co_io_inputs_codewords_2),
    .io_inputs_codewords_3(co_io_inputs_codewords_3),
    .io_inputs_codewords_4(co_io_inputs_codewords_4),
    .io_inputs_codewords_5(co_io_inputs_codewords_5),
    .io_inputs_codewords_6(co_io_inputs_codewords_6),
    .io_inputs_codewords_7(co_io_inputs_codewords_7),
    .io_inputs_codewords_8(co_io_inputs_codewords_8),
    .io_inputs_codewords_9(co_io_inputs_codewords_9),
    .io_inputs_codewords_10(co_io_inputs_codewords_10),
    .io_inputs_codewords_11(co_io_inputs_codewords_11),
    .io_inputs_codewords_12(co_io_inputs_codewords_12),
    .io_inputs_codewords_13(co_io_inputs_codewords_13),
    .io_inputs_codewords_14(co_io_inputs_codewords_14),
    .io_inputs_codewords_15(co_io_inputs_codewords_15),
    .io_inputs_codewords_16(co_io_inputs_codewords_16),
    .io_inputs_codewords_17(co_io_inputs_codewords_17),
    .io_inputs_codewords_18(co_io_inputs_codewords_18),
    .io_inputs_codewords_19(co_io_inputs_codewords_19),
    .io_inputs_codewords_20(co_io_inputs_codewords_20),
    .io_inputs_codewords_21(co_io_inputs_codewords_21),
    .io_inputs_codewords_22(co_io_inputs_codewords_22),
    .io_inputs_codewords_23(co_io_inputs_codewords_23),
    .io_inputs_codewords_24(co_io_inputs_codewords_24),
    .io_inputs_codewords_25(co_io_inputs_codewords_25),
    .io_inputs_codewords_26(co_io_inputs_codewords_26),
    .io_inputs_codewords_27(co_io_inputs_codewords_27),
    .io_inputs_codewords_28(co_io_inputs_codewords_28),
    .io_inputs_codewords_29(co_io_inputs_codewords_29),
    .io_inputs_codewords_30(co_io_inputs_codewords_30),
    .io_inputs_codewords_31(co_io_inputs_codewords_31),
    .io_inputs_codewords_32(co_io_inputs_codewords_32),
    .io_inputs_codewords_33(co_io_inputs_codewords_33),
    .io_inputs_codewords_34(co_io_inputs_codewords_34),
    .io_inputs_codewords_35(co_io_inputs_codewords_35),
    .io_inputs_codewords_36(co_io_inputs_codewords_36),
    .io_inputs_codewords_37(co_io_inputs_codewords_37),
    .io_inputs_codewords_38(co_io_inputs_codewords_38),
    .io_inputs_codewords_39(co_io_inputs_codewords_39),
    .io_inputs_codewords_40(co_io_inputs_codewords_40),
    .io_inputs_codewords_41(co_io_inputs_codewords_41),
    .io_inputs_codewords_42(co_io_inputs_codewords_42),
    .io_inputs_codewords_43(co_io_inputs_codewords_43),
    .io_inputs_codewords_44(co_io_inputs_codewords_44),
    .io_inputs_codewords_45(co_io_inputs_codewords_45),
    .io_inputs_codewords_46(co_io_inputs_codewords_46),
    .io_inputs_codewords_47(co_io_inputs_codewords_47),
    .io_inputs_codewords_48(co_io_inputs_codewords_48),
    .io_inputs_codewords_49(co_io_inputs_codewords_49),
    .io_inputs_codewords_50(co_io_inputs_codewords_50),
    .io_inputs_codewords_51(co_io_inputs_codewords_51),
    .io_inputs_codewords_52(co_io_inputs_codewords_52),
    .io_inputs_codewords_53(co_io_inputs_codewords_53),
    .io_inputs_codewords_54(co_io_inputs_codewords_54),
    .io_inputs_codewords_55(co_io_inputs_codewords_55),
    .io_inputs_codewords_56(co_io_inputs_codewords_56),
    .io_inputs_codewords_57(co_io_inputs_codewords_57),
    .io_inputs_codewords_58(co_io_inputs_codewords_58),
    .io_inputs_codewords_59(co_io_inputs_codewords_59),
    .io_inputs_codewords_60(co_io_inputs_codewords_60),
    .io_inputs_codewords_61(co_io_inputs_codewords_61),
    .io_inputs_codewords_62(co_io_inputs_codewords_62),
    .io_inputs_codewords_63(co_io_inputs_codewords_63),
    .io_inputs_codewords_64(co_io_inputs_codewords_64),
    .io_inputs_codewords_65(co_io_inputs_codewords_65),
    .io_inputs_codewords_66(co_io_inputs_codewords_66),
    .io_inputs_codewords_67(co_io_inputs_codewords_67),
    .io_inputs_codewords_68(co_io_inputs_codewords_68),
    .io_inputs_codewords_69(co_io_inputs_codewords_69),
    .io_inputs_codewords_70(co_io_inputs_codewords_70),
    .io_inputs_codewords_71(co_io_inputs_codewords_71),
    .io_inputs_codewords_72(co_io_inputs_codewords_72),
    .io_inputs_codewords_73(co_io_inputs_codewords_73),
    .io_inputs_codewords_74(co_io_inputs_codewords_74),
    .io_inputs_codewords_75(co_io_inputs_codewords_75),
    .io_inputs_codewords_76(co_io_inputs_codewords_76),
    .io_inputs_codewords_77(co_io_inputs_codewords_77),
    .io_inputs_codewords_78(co_io_inputs_codewords_78),
    .io_inputs_codewords_79(co_io_inputs_codewords_79),
    .io_inputs_codewords_80(co_io_inputs_codewords_80),
    .io_inputs_codewords_81(co_io_inputs_codewords_81),
    .io_inputs_codewords_82(co_io_inputs_codewords_82),
    .io_inputs_codewords_83(co_io_inputs_codewords_83),
    .io_inputs_codewords_84(co_io_inputs_codewords_84),
    .io_inputs_codewords_85(co_io_inputs_codewords_85),
    .io_inputs_codewords_86(co_io_inputs_codewords_86),
    .io_inputs_codewords_87(co_io_inputs_codewords_87),
    .io_inputs_codewords_88(co_io_inputs_codewords_88),
    .io_inputs_codewords_89(co_io_inputs_codewords_89),
    .io_inputs_codewords_90(co_io_inputs_codewords_90),
    .io_inputs_codewords_91(co_io_inputs_codewords_91),
    .io_inputs_codewords_92(co_io_inputs_codewords_92),
    .io_inputs_codewords_93(co_io_inputs_codewords_93),
    .io_inputs_codewords_94(co_io_inputs_codewords_94),
    .io_inputs_codewords_95(co_io_inputs_codewords_95),
    .io_inputs_codewords_96(co_io_inputs_codewords_96),
    .io_inputs_codewords_97(co_io_inputs_codewords_97),
    .io_inputs_codewords_98(co_io_inputs_codewords_98),
    .io_inputs_codewords_99(co_io_inputs_codewords_99),
    .io_inputs_codewords_100(co_io_inputs_codewords_100),
    .io_inputs_codewords_101(co_io_inputs_codewords_101),
    .io_inputs_codewords_102(co_io_inputs_codewords_102),
    .io_inputs_codewords_103(co_io_inputs_codewords_103),
    .io_inputs_codewords_104(co_io_inputs_codewords_104),
    .io_inputs_codewords_105(co_io_inputs_codewords_105),
    .io_inputs_codewords_106(co_io_inputs_codewords_106),
    .io_inputs_codewords_107(co_io_inputs_codewords_107),
    .io_inputs_codewords_108(co_io_inputs_codewords_108),
    .io_inputs_codewords_109(co_io_inputs_codewords_109),
    .io_inputs_codewords_110(co_io_inputs_codewords_110),
    .io_inputs_codewords_111(co_io_inputs_codewords_111),
    .io_inputs_codewords_112(co_io_inputs_codewords_112),
    .io_inputs_codewords_113(co_io_inputs_codewords_113),
    .io_inputs_codewords_114(co_io_inputs_codewords_114),
    .io_inputs_codewords_115(co_io_inputs_codewords_115),
    .io_inputs_codewords_116(co_io_inputs_codewords_116),
    .io_inputs_codewords_117(co_io_inputs_codewords_117),
    .io_inputs_codewords_118(co_io_inputs_codewords_118),
    .io_inputs_codewords_119(co_io_inputs_codewords_119),
    .io_inputs_codewords_120(co_io_inputs_codewords_120),
    .io_inputs_codewords_121(co_io_inputs_codewords_121),
    .io_inputs_codewords_122(co_io_inputs_codewords_122),
    .io_inputs_codewords_123(co_io_inputs_codewords_123),
    .io_inputs_codewords_124(co_io_inputs_codewords_124),
    .io_inputs_codewords_125(co_io_inputs_codewords_125),
    .io_inputs_codewords_126(co_io_inputs_codewords_126),
    .io_inputs_codewords_127(co_io_inputs_codewords_127),
    .io_inputs_codewords_128(co_io_inputs_codewords_128),
    .io_inputs_codewords_129(co_io_inputs_codewords_129),
    .io_inputs_codewords_130(co_io_inputs_codewords_130),
    .io_inputs_codewords_131(co_io_inputs_codewords_131),
    .io_inputs_codewords_132(co_io_inputs_codewords_132),
    .io_inputs_codewords_133(co_io_inputs_codewords_133),
    .io_inputs_codewords_134(co_io_inputs_codewords_134),
    .io_inputs_codewords_135(co_io_inputs_codewords_135),
    .io_inputs_codewords_136(co_io_inputs_codewords_136),
    .io_inputs_codewords_137(co_io_inputs_codewords_137),
    .io_inputs_codewords_138(co_io_inputs_codewords_138),
    .io_inputs_codewords_139(co_io_inputs_codewords_139),
    .io_inputs_codewords_140(co_io_inputs_codewords_140),
    .io_inputs_codewords_141(co_io_inputs_codewords_141),
    .io_inputs_codewords_142(co_io_inputs_codewords_142),
    .io_inputs_codewords_143(co_io_inputs_codewords_143),
    .io_inputs_codewords_144(co_io_inputs_codewords_144),
    .io_inputs_codewords_145(co_io_inputs_codewords_145),
    .io_inputs_codewords_146(co_io_inputs_codewords_146),
    .io_inputs_codewords_147(co_io_inputs_codewords_147),
    .io_inputs_codewords_148(co_io_inputs_codewords_148),
    .io_inputs_codewords_149(co_io_inputs_codewords_149),
    .io_inputs_codewords_150(co_io_inputs_codewords_150),
    .io_inputs_codewords_151(co_io_inputs_codewords_151),
    .io_inputs_codewords_152(co_io_inputs_codewords_152),
    .io_inputs_codewords_153(co_io_inputs_codewords_153),
    .io_inputs_codewords_154(co_io_inputs_codewords_154),
    .io_inputs_codewords_155(co_io_inputs_codewords_155),
    .io_inputs_codewords_156(co_io_inputs_codewords_156),
    .io_inputs_codewords_157(co_io_inputs_codewords_157),
    .io_inputs_codewords_158(co_io_inputs_codewords_158),
    .io_inputs_codewords_159(co_io_inputs_codewords_159),
    .io_inputs_codewords_160(co_io_inputs_codewords_160),
    .io_inputs_codewords_161(co_io_inputs_codewords_161),
    .io_inputs_codewords_162(co_io_inputs_codewords_162),
    .io_inputs_codewords_163(co_io_inputs_codewords_163),
    .io_inputs_codewords_164(co_io_inputs_codewords_164),
    .io_inputs_codewords_165(co_io_inputs_codewords_165),
    .io_inputs_codewords_166(co_io_inputs_codewords_166),
    .io_inputs_codewords_167(co_io_inputs_codewords_167),
    .io_inputs_codewords_168(co_io_inputs_codewords_168),
    .io_inputs_codewords_169(co_io_inputs_codewords_169),
    .io_inputs_codewords_170(co_io_inputs_codewords_170),
    .io_inputs_codewords_171(co_io_inputs_codewords_171),
    .io_inputs_codewords_172(co_io_inputs_codewords_172),
    .io_inputs_codewords_173(co_io_inputs_codewords_173),
    .io_inputs_codewords_174(co_io_inputs_codewords_174),
    .io_inputs_codewords_175(co_io_inputs_codewords_175),
    .io_inputs_codewords_176(co_io_inputs_codewords_176),
    .io_inputs_codewords_177(co_io_inputs_codewords_177),
    .io_inputs_codewords_178(co_io_inputs_codewords_178),
    .io_inputs_codewords_179(co_io_inputs_codewords_179),
    .io_inputs_codewords_180(co_io_inputs_codewords_180),
    .io_inputs_codewords_181(co_io_inputs_codewords_181),
    .io_inputs_codewords_182(co_io_inputs_codewords_182),
    .io_inputs_codewords_183(co_io_inputs_codewords_183),
    .io_inputs_codewords_184(co_io_inputs_codewords_184),
    .io_inputs_codewords_185(co_io_inputs_codewords_185),
    .io_inputs_codewords_186(co_io_inputs_codewords_186),
    .io_inputs_codewords_187(co_io_inputs_codewords_187),
    .io_inputs_codewords_188(co_io_inputs_codewords_188),
    .io_inputs_codewords_189(co_io_inputs_codewords_189),
    .io_inputs_codewords_190(co_io_inputs_codewords_190),
    .io_inputs_codewords_191(co_io_inputs_codewords_191),
    .io_inputs_codewords_192(co_io_inputs_codewords_192),
    .io_inputs_codewords_193(co_io_inputs_codewords_193),
    .io_inputs_codewords_194(co_io_inputs_codewords_194),
    .io_inputs_codewords_195(co_io_inputs_codewords_195),
    .io_inputs_codewords_196(co_io_inputs_codewords_196),
    .io_inputs_codewords_197(co_io_inputs_codewords_197),
    .io_inputs_codewords_198(co_io_inputs_codewords_198),
    .io_inputs_codewords_199(co_io_inputs_codewords_199),
    .io_inputs_codewords_200(co_io_inputs_codewords_200),
    .io_inputs_codewords_201(co_io_inputs_codewords_201),
    .io_inputs_codewords_202(co_io_inputs_codewords_202),
    .io_inputs_codewords_203(co_io_inputs_codewords_203),
    .io_inputs_codewords_204(co_io_inputs_codewords_204),
    .io_inputs_codewords_205(co_io_inputs_codewords_205),
    .io_inputs_codewords_206(co_io_inputs_codewords_206),
    .io_inputs_codewords_207(co_io_inputs_codewords_207),
    .io_inputs_codewords_208(co_io_inputs_codewords_208),
    .io_inputs_codewords_209(co_io_inputs_codewords_209),
    .io_inputs_codewords_210(co_io_inputs_codewords_210),
    .io_inputs_codewords_211(co_io_inputs_codewords_211),
    .io_inputs_codewords_212(co_io_inputs_codewords_212),
    .io_inputs_codewords_213(co_io_inputs_codewords_213),
    .io_inputs_codewords_214(co_io_inputs_codewords_214),
    .io_inputs_codewords_215(co_io_inputs_codewords_215),
    .io_inputs_codewords_216(co_io_inputs_codewords_216),
    .io_inputs_codewords_217(co_io_inputs_codewords_217),
    .io_inputs_codewords_218(co_io_inputs_codewords_218),
    .io_inputs_codewords_219(co_io_inputs_codewords_219),
    .io_inputs_codewords_220(co_io_inputs_codewords_220),
    .io_inputs_codewords_221(co_io_inputs_codewords_221),
    .io_inputs_codewords_222(co_io_inputs_codewords_222),
    .io_inputs_codewords_223(co_io_inputs_codewords_223),
    .io_inputs_codewords_224(co_io_inputs_codewords_224),
    .io_inputs_codewords_225(co_io_inputs_codewords_225),
    .io_inputs_codewords_226(co_io_inputs_codewords_226),
    .io_inputs_codewords_227(co_io_inputs_codewords_227),
    .io_inputs_codewords_228(co_io_inputs_codewords_228),
    .io_inputs_codewords_229(co_io_inputs_codewords_229),
    .io_inputs_codewords_230(co_io_inputs_codewords_230),
    .io_inputs_codewords_231(co_io_inputs_codewords_231),
    .io_inputs_codewords_232(co_io_inputs_codewords_232),
    .io_inputs_codewords_233(co_io_inputs_codewords_233),
    .io_inputs_codewords_234(co_io_inputs_codewords_234),
    .io_inputs_codewords_235(co_io_inputs_codewords_235),
    .io_inputs_codewords_236(co_io_inputs_codewords_236),
    .io_inputs_codewords_237(co_io_inputs_codewords_237),
    .io_inputs_codewords_238(co_io_inputs_codewords_238),
    .io_inputs_codewords_239(co_io_inputs_codewords_239),
    .io_inputs_codewords_240(co_io_inputs_codewords_240),
    .io_inputs_codewords_241(co_io_inputs_codewords_241),
    .io_inputs_codewords_242(co_io_inputs_codewords_242),
    .io_inputs_codewords_243(co_io_inputs_codewords_243),
    .io_inputs_codewords_244(co_io_inputs_codewords_244),
    .io_inputs_codewords_245(co_io_inputs_codewords_245),
    .io_inputs_codewords_246(co_io_inputs_codewords_246),
    .io_inputs_codewords_247(co_io_inputs_codewords_247),
    .io_inputs_codewords_248(co_io_inputs_codewords_248),
    .io_inputs_codewords_249(co_io_inputs_codewords_249),
    .io_inputs_codewords_250(co_io_inputs_codewords_250),
    .io_inputs_codewords_251(co_io_inputs_codewords_251),
    .io_inputs_codewords_252(co_io_inputs_codewords_252),
    .io_inputs_codewords_253(co_io_inputs_codewords_253),
    .io_inputs_codewords_254(co_io_inputs_codewords_254),
    .io_inputs_codewords_255(co_io_inputs_codewords_255),
    .io_inputs_lengths_0(co_io_inputs_lengths_0),
    .io_inputs_lengths_1(co_io_inputs_lengths_1),
    .io_inputs_lengths_2(co_io_inputs_lengths_2),
    .io_inputs_lengths_3(co_io_inputs_lengths_3),
    .io_inputs_lengths_4(co_io_inputs_lengths_4),
    .io_inputs_lengths_5(co_io_inputs_lengths_5),
    .io_inputs_lengths_6(co_io_inputs_lengths_6),
    .io_inputs_lengths_7(co_io_inputs_lengths_7),
    .io_inputs_lengths_8(co_io_inputs_lengths_8),
    .io_inputs_lengths_9(co_io_inputs_lengths_9),
    .io_inputs_lengths_10(co_io_inputs_lengths_10),
    .io_inputs_lengths_11(co_io_inputs_lengths_11),
    .io_inputs_lengths_12(co_io_inputs_lengths_12),
    .io_inputs_lengths_13(co_io_inputs_lengths_13),
    .io_inputs_lengths_14(co_io_inputs_lengths_14),
    .io_inputs_lengths_15(co_io_inputs_lengths_15),
    .io_inputs_lengths_16(co_io_inputs_lengths_16),
    .io_inputs_lengths_17(co_io_inputs_lengths_17),
    .io_inputs_lengths_18(co_io_inputs_lengths_18),
    .io_inputs_lengths_19(co_io_inputs_lengths_19),
    .io_inputs_lengths_20(co_io_inputs_lengths_20),
    .io_inputs_lengths_21(co_io_inputs_lengths_21),
    .io_inputs_lengths_22(co_io_inputs_lengths_22),
    .io_inputs_lengths_23(co_io_inputs_lengths_23),
    .io_inputs_lengths_24(co_io_inputs_lengths_24),
    .io_inputs_lengths_25(co_io_inputs_lengths_25),
    .io_inputs_lengths_26(co_io_inputs_lengths_26),
    .io_inputs_lengths_27(co_io_inputs_lengths_27),
    .io_inputs_lengths_28(co_io_inputs_lengths_28),
    .io_inputs_lengths_29(co_io_inputs_lengths_29),
    .io_inputs_lengths_30(co_io_inputs_lengths_30),
    .io_inputs_lengths_31(co_io_inputs_lengths_31),
    .io_inputs_lengths_32(co_io_inputs_lengths_32),
    .io_inputs_lengths_33(co_io_inputs_lengths_33),
    .io_inputs_lengths_34(co_io_inputs_lengths_34),
    .io_inputs_lengths_35(co_io_inputs_lengths_35),
    .io_inputs_lengths_36(co_io_inputs_lengths_36),
    .io_inputs_lengths_37(co_io_inputs_lengths_37),
    .io_inputs_lengths_38(co_io_inputs_lengths_38),
    .io_inputs_lengths_39(co_io_inputs_lengths_39),
    .io_inputs_lengths_40(co_io_inputs_lengths_40),
    .io_inputs_lengths_41(co_io_inputs_lengths_41),
    .io_inputs_lengths_42(co_io_inputs_lengths_42),
    .io_inputs_lengths_43(co_io_inputs_lengths_43),
    .io_inputs_lengths_44(co_io_inputs_lengths_44),
    .io_inputs_lengths_45(co_io_inputs_lengths_45),
    .io_inputs_lengths_46(co_io_inputs_lengths_46),
    .io_inputs_lengths_47(co_io_inputs_lengths_47),
    .io_inputs_lengths_48(co_io_inputs_lengths_48),
    .io_inputs_lengths_49(co_io_inputs_lengths_49),
    .io_inputs_lengths_50(co_io_inputs_lengths_50),
    .io_inputs_lengths_51(co_io_inputs_lengths_51),
    .io_inputs_lengths_52(co_io_inputs_lengths_52),
    .io_inputs_lengths_53(co_io_inputs_lengths_53),
    .io_inputs_lengths_54(co_io_inputs_lengths_54),
    .io_inputs_lengths_55(co_io_inputs_lengths_55),
    .io_inputs_lengths_56(co_io_inputs_lengths_56),
    .io_inputs_lengths_57(co_io_inputs_lengths_57),
    .io_inputs_lengths_58(co_io_inputs_lengths_58),
    .io_inputs_lengths_59(co_io_inputs_lengths_59),
    .io_inputs_lengths_60(co_io_inputs_lengths_60),
    .io_inputs_lengths_61(co_io_inputs_lengths_61),
    .io_inputs_lengths_62(co_io_inputs_lengths_62),
    .io_inputs_lengths_63(co_io_inputs_lengths_63),
    .io_inputs_lengths_64(co_io_inputs_lengths_64),
    .io_inputs_lengths_65(co_io_inputs_lengths_65),
    .io_inputs_lengths_66(co_io_inputs_lengths_66),
    .io_inputs_lengths_67(co_io_inputs_lengths_67),
    .io_inputs_lengths_68(co_io_inputs_lengths_68),
    .io_inputs_lengths_69(co_io_inputs_lengths_69),
    .io_inputs_lengths_70(co_io_inputs_lengths_70),
    .io_inputs_lengths_71(co_io_inputs_lengths_71),
    .io_inputs_lengths_72(co_io_inputs_lengths_72),
    .io_inputs_lengths_73(co_io_inputs_lengths_73),
    .io_inputs_lengths_74(co_io_inputs_lengths_74),
    .io_inputs_lengths_75(co_io_inputs_lengths_75),
    .io_inputs_lengths_76(co_io_inputs_lengths_76),
    .io_inputs_lengths_77(co_io_inputs_lengths_77),
    .io_inputs_lengths_78(co_io_inputs_lengths_78),
    .io_inputs_lengths_79(co_io_inputs_lengths_79),
    .io_inputs_lengths_80(co_io_inputs_lengths_80),
    .io_inputs_lengths_81(co_io_inputs_lengths_81),
    .io_inputs_lengths_82(co_io_inputs_lengths_82),
    .io_inputs_lengths_83(co_io_inputs_lengths_83),
    .io_inputs_lengths_84(co_io_inputs_lengths_84),
    .io_inputs_lengths_85(co_io_inputs_lengths_85),
    .io_inputs_lengths_86(co_io_inputs_lengths_86),
    .io_inputs_lengths_87(co_io_inputs_lengths_87),
    .io_inputs_lengths_88(co_io_inputs_lengths_88),
    .io_inputs_lengths_89(co_io_inputs_lengths_89),
    .io_inputs_lengths_90(co_io_inputs_lengths_90),
    .io_inputs_lengths_91(co_io_inputs_lengths_91),
    .io_inputs_lengths_92(co_io_inputs_lengths_92),
    .io_inputs_lengths_93(co_io_inputs_lengths_93),
    .io_inputs_lengths_94(co_io_inputs_lengths_94),
    .io_inputs_lengths_95(co_io_inputs_lengths_95),
    .io_inputs_lengths_96(co_io_inputs_lengths_96),
    .io_inputs_lengths_97(co_io_inputs_lengths_97),
    .io_inputs_lengths_98(co_io_inputs_lengths_98),
    .io_inputs_lengths_99(co_io_inputs_lengths_99),
    .io_inputs_lengths_100(co_io_inputs_lengths_100),
    .io_inputs_lengths_101(co_io_inputs_lengths_101),
    .io_inputs_lengths_102(co_io_inputs_lengths_102),
    .io_inputs_lengths_103(co_io_inputs_lengths_103),
    .io_inputs_lengths_104(co_io_inputs_lengths_104),
    .io_inputs_lengths_105(co_io_inputs_lengths_105),
    .io_inputs_lengths_106(co_io_inputs_lengths_106),
    .io_inputs_lengths_107(co_io_inputs_lengths_107),
    .io_inputs_lengths_108(co_io_inputs_lengths_108),
    .io_inputs_lengths_109(co_io_inputs_lengths_109),
    .io_inputs_lengths_110(co_io_inputs_lengths_110),
    .io_inputs_lengths_111(co_io_inputs_lengths_111),
    .io_inputs_lengths_112(co_io_inputs_lengths_112),
    .io_inputs_lengths_113(co_io_inputs_lengths_113),
    .io_inputs_lengths_114(co_io_inputs_lengths_114),
    .io_inputs_lengths_115(co_io_inputs_lengths_115),
    .io_inputs_lengths_116(co_io_inputs_lengths_116),
    .io_inputs_lengths_117(co_io_inputs_lengths_117),
    .io_inputs_lengths_118(co_io_inputs_lengths_118),
    .io_inputs_lengths_119(co_io_inputs_lengths_119),
    .io_inputs_lengths_120(co_io_inputs_lengths_120),
    .io_inputs_lengths_121(co_io_inputs_lengths_121),
    .io_inputs_lengths_122(co_io_inputs_lengths_122),
    .io_inputs_lengths_123(co_io_inputs_lengths_123),
    .io_inputs_lengths_124(co_io_inputs_lengths_124),
    .io_inputs_lengths_125(co_io_inputs_lengths_125),
    .io_inputs_lengths_126(co_io_inputs_lengths_126),
    .io_inputs_lengths_127(co_io_inputs_lengths_127),
    .io_inputs_lengths_128(co_io_inputs_lengths_128),
    .io_inputs_lengths_129(co_io_inputs_lengths_129),
    .io_inputs_lengths_130(co_io_inputs_lengths_130),
    .io_inputs_lengths_131(co_io_inputs_lengths_131),
    .io_inputs_lengths_132(co_io_inputs_lengths_132),
    .io_inputs_lengths_133(co_io_inputs_lengths_133),
    .io_inputs_lengths_134(co_io_inputs_lengths_134),
    .io_inputs_lengths_135(co_io_inputs_lengths_135),
    .io_inputs_lengths_136(co_io_inputs_lengths_136),
    .io_inputs_lengths_137(co_io_inputs_lengths_137),
    .io_inputs_lengths_138(co_io_inputs_lengths_138),
    .io_inputs_lengths_139(co_io_inputs_lengths_139),
    .io_inputs_lengths_140(co_io_inputs_lengths_140),
    .io_inputs_lengths_141(co_io_inputs_lengths_141),
    .io_inputs_lengths_142(co_io_inputs_lengths_142),
    .io_inputs_lengths_143(co_io_inputs_lengths_143),
    .io_inputs_lengths_144(co_io_inputs_lengths_144),
    .io_inputs_lengths_145(co_io_inputs_lengths_145),
    .io_inputs_lengths_146(co_io_inputs_lengths_146),
    .io_inputs_lengths_147(co_io_inputs_lengths_147),
    .io_inputs_lengths_148(co_io_inputs_lengths_148),
    .io_inputs_lengths_149(co_io_inputs_lengths_149),
    .io_inputs_lengths_150(co_io_inputs_lengths_150),
    .io_inputs_lengths_151(co_io_inputs_lengths_151),
    .io_inputs_lengths_152(co_io_inputs_lengths_152),
    .io_inputs_lengths_153(co_io_inputs_lengths_153),
    .io_inputs_lengths_154(co_io_inputs_lengths_154),
    .io_inputs_lengths_155(co_io_inputs_lengths_155),
    .io_inputs_lengths_156(co_io_inputs_lengths_156),
    .io_inputs_lengths_157(co_io_inputs_lengths_157),
    .io_inputs_lengths_158(co_io_inputs_lengths_158),
    .io_inputs_lengths_159(co_io_inputs_lengths_159),
    .io_inputs_lengths_160(co_io_inputs_lengths_160),
    .io_inputs_lengths_161(co_io_inputs_lengths_161),
    .io_inputs_lengths_162(co_io_inputs_lengths_162),
    .io_inputs_lengths_163(co_io_inputs_lengths_163),
    .io_inputs_lengths_164(co_io_inputs_lengths_164),
    .io_inputs_lengths_165(co_io_inputs_lengths_165),
    .io_inputs_lengths_166(co_io_inputs_lengths_166),
    .io_inputs_lengths_167(co_io_inputs_lengths_167),
    .io_inputs_lengths_168(co_io_inputs_lengths_168),
    .io_inputs_lengths_169(co_io_inputs_lengths_169),
    .io_inputs_lengths_170(co_io_inputs_lengths_170),
    .io_inputs_lengths_171(co_io_inputs_lengths_171),
    .io_inputs_lengths_172(co_io_inputs_lengths_172),
    .io_inputs_lengths_173(co_io_inputs_lengths_173),
    .io_inputs_lengths_174(co_io_inputs_lengths_174),
    .io_inputs_lengths_175(co_io_inputs_lengths_175),
    .io_inputs_lengths_176(co_io_inputs_lengths_176),
    .io_inputs_lengths_177(co_io_inputs_lengths_177),
    .io_inputs_lengths_178(co_io_inputs_lengths_178),
    .io_inputs_lengths_179(co_io_inputs_lengths_179),
    .io_inputs_lengths_180(co_io_inputs_lengths_180),
    .io_inputs_lengths_181(co_io_inputs_lengths_181),
    .io_inputs_lengths_182(co_io_inputs_lengths_182),
    .io_inputs_lengths_183(co_io_inputs_lengths_183),
    .io_inputs_lengths_184(co_io_inputs_lengths_184),
    .io_inputs_lengths_185(co_io_inputs_lengths_185),
    .io_inputs_lengths_186(co_io_inputs_lengths_186),
    .io_inputs_lengths_187(co_io_inputs_lengths_187),
    .io_inputs_lengths_188(co_io_inputs_lengths_188),
    .io_inputs_lengths_189(co_io_inputs_lengths_189),
    .io_inputs_lengths_190(co_io_inputs_lengths_190),
    .io_inputs_lengths_191(co_io_inputs_lengths_191),
    .io_inputs_lengths_192(co_io_inputs_lengths_192),
    .io_inputs_lengths_193(co_io_inputs_lengths_193),
    .io_inputs_lengths_194(co_io_inputs_lengths_194),
    .io_inputs_lengths_195(co_io_inputs_lengths_195),
    .io_inputs_lengths_196(co_io_inputs_lengths_196),
    .io_inputs_lengths_197(co_io_inputs_lengths_197),
    .io_inputs_lengths_198(co_io_inputs_lengths_198),
    .io_inputs_lengths_199(co_io_inputs_lengths_199),
    .io_inputs_lengths_200(co_io_inputs_lengths_200),
    .io_inputs_lengths_201(co_io_inputs_lengths_201),
    .io_inputs_lengths_202(co_io_inputs_lengths_202),
    .io_inputs_lengths_203(co_io_inputs_lengths_203),
    .io_inputs_lengths_204(co_io_inputs_lengths_204),
    .io_inputs_lengths_205(co_io_inputs_lengths_205),
    .io_inputs_lengths_206(co_io_inputs_lengths_206),
    .io_inputs_lengths_207(co_io_inputs_lengths_207),
    .io_inputs_lengths_208(co_io_inputs_lengths_208),
    .io_inputs_lengths_209(co_io_inputs_lengths_209),
    .io_inputs_lengths_210(co_io_inputs_lengths_210),
    .io_inputs_lengths_211(co_io_inputs_lengths_211),
    .io_inputs_lengths_212(co_io_inputs_lengths_212),
    .io_inputs_lengths_213(co_io_inputs_lengths_213),
    .io_inputs_lengths_214(co_io_inputs_lengths_214),
    .io_inputs_lengths_215(co_io_inputs_lengths_215),
    .io_inputs_lengths_216(co_io_inputs_lengths_216),
    .io_inputs_lengths_217(co_io_inputs_lengths_217),
    .io_inputs_lengths_218(co_io_inputs_lengths_218),
    .io_inputs_lengths_219(co_io_inputs_lengths_219),
    .io_inputs_lengths_220(co_io_inputs_lengths_220),
    .io_inputs_lengths_221(co_io_inputs_lengths_221),
    .io_inputs_lengths_222(co_io_inputs_lengths_222),
    .io_inputs_lengths_223(co_io_inputs_lengths_223),
    .io_inputs_lengths_224(co_io_inputs_lengths_224),
    .io_inputs_lengths_225(co_io_inputs_lengths_225),
    .io_inputs_lengths_226(co_io_inputs_lengths_226),
    .io_inputs_lengths_227(co_io_inputs_lengths_227),
    .io_inputs_lengths_228(co_io_inputs_lengths_228),
    .io_inputs_lengths_229(co_io_inputs_lengths_229),
    .io_inputs_lengths_230(co_io_inputs_lengths_230),
    .io_inputs_lengths_231(co_io_inputs_lengths_231),
    .io_inputs_lengths_232(co_io_inputs_lengths_232),
    .io_inputs_lengths_233(co_io_inputs_lengths_233),
    .io_inputs_lengths_234(co_io_inputs_lengths_234),
    .io_inputs_lengths_235(co_io_inputs_lengths_235),
    .io_inputs_lengths_236(co_io_inputs_lengths_236),
    .io_inputs_lengths_237(co_io_inputs_lengths_237),
    .io_inputs_lengths_238(co_io_inputs_lengths_238),
    .io_inputs_lengths_239(co_io_inputs_lengths_239),
    .io_inputs_lengths_240(co_io_inputs_lengths_240),
    .io_inputs_lengths_241(co_io_inputs_lengths_241),
    .io_inputs_lengths_242(co_io_inputs_lengths_242),
    .io_inputs_lengths_243(co_io_inputs_lengths_243),
    .io_inputs_lengths_244(co_io_inputs_lengths_244),
    .io_inputs_lengths_245(co_io_inputs_lengths_245),
    .io_inputs_lengths_246(co_io_inputs_lengths_246),
    .io_inputs_lengths_247(co_io_inputs_lengths_247),
    .io_inputs_lengths_248(co_io_inputs_lengths_248),
    .io_inputs_lengths_249(co_io_inputs_lengths_249),
    .io_inputs_lengths_250(co_io_inputs_lengths_250),
    .io_inputs_lengths_251(co_io_inputs_lengths_251),
    .io_inputs_lengths_252(co_io_inputs_lengths_252),
    .io_inputs_lengths_253(co_io_inputs_lengths_253),
    .io_inputs_lengths_254(co_io_inputs_lengths_254),
    .io_inputs_lengths_255(co_io_inputs_lengths_255),
    .io_inputs_charactersOut_0(co_io_inputs_charactersOut_0),
    .io_inputs_charactersOut_1(co_io_inputs_charactersOut_1),
    .io_inputs_charactersOut_2(co_io_inputs_charactersOut_2),
    .io_inputs_charactersOut_3(co_io_inputs_charactersOut_3),
    .io_inputs_charactersOut_4(co_io_inputs_charactersOut_4),
    .io_inputs_charactersOut_5(co_io_inputs_charactersOut_5),
    .io_inputs_charactersOut_6(co_io_inputs_charactersOut_6),
    .io_inputs_charactersOut_7(co_io_inputs_charactersOut_7),
    .io_inputs_charactersOut_8(co_io_inputs_charactersOut_8),
    .io_inputs_charactersOut_9(co_io_inputs_charactersOut_9),
    .io_inputs_charactersOut_10(co_io_inputs_charactersOut_10),
    .io_inputs_charactersOut_11(co_io_inputs_charactersOut_11),
    .io_inputs_charactersOut_12(co_io_inputs_charactersOut_12),
    .io_inputs_charactersOut_13(co_io_inputs_charactersOut_13),
    .io_inputs_charactersOut_14(co_io_inputs_charactersOut_14),
    .io_inputs_charactersOut_15(co_io_inputs_charactersOut_15),
    .io_inputs_charactersOut_16(co_io_inputs_charactersOut_16),
    .io_inputs_charactersOut_17(co_io_inputs_charactersOut_17),
    .io_inputs_charactersOut_18(co_io_inputs_charactersOut_18),
    .io_inputs_charactersOut_19(co_io_inputs_charactersOut_19),
    .io_inputs_charactersOut_20(co_io_inputs_charactersOut_20),
    .io_inputs_charactersOut_21(co_io_inputs_charactersOut_21),
    .io_inputs_charactersOut_22(co_io_inputs_charactersOut_22),
    .io_inputs_charactersOut_23(co_io_inputs_charactersOut_23),
    .io_inputs_charactersOut_24(co_io_inputs_charactersOut_24),
    .io_inputs_charactersOut_25(co_io_inputs_charactersOut_25),
    .io_inputs_charactersOut_26(co_io_inputs_charactersOut_26),
    .io_inputs_charactersOut_27(co_io_inputs_charactersOut_27),
    .io_inputs_charactersOut_28(co_io_inputs_charactersOut_28),
    .io_inputs_charactersOut_29(co_io_inputs_charactersOut_29),
    .io_inputs_charactersOut_30(co_io_inputs_charactersOut_30),
    .io_inputs_charactersOut_31(co_io_inputs_charactersOut_31),
    .io_inputs_nodes(co_io_inputs_nodes),
    .io_inputs_escapeCharacterLength(co_io_inputs_escapeCharacterLength),
    .io_inputs_escapeCodeword(co_io_inputs_escapeCodeword),
    .io_outputs_0_dataOut(co_io_outputs_0_dataOut),
    .io_outputs_0_dataLength(co_io_outputs_0_dataLength),
    .io_outputs_0_valid(co_io_outputs_0_valid),
    .io_outputs_0_ready(co_io_outputs_0_ready),
    .io_finished(co_io_finished)
  );
  assign io_characterFrequencyInputs_currentByteOut = cfm_io_input_currentByteOut; // @[topLevel.scala 93:31]
  assign io_characterFrequencyInputs_ready = cfm_io_input_ready; // @[topLevel.scala 93:31]
  assign io_compressionInputs_0_currentByteOut = co_io_dataIn_0_currentByteOut; // @[topLevel.scala 95:33]
  assign io_compressionInputs_0_ready = co_io_dataIn_0_ready; // @[topLevel.scala 95:33]
  assign io_outputs_0_dataOut = co_io_outputs_0_dataOut; // @[topLevel.scala 103:14]
  assign io_outputs_0_dataLength = co_io_outputs_0_dataLength; // @[topLevel.scala 103:14]
  assign io_outputs_0_valid = co_io_outputs_0_valid; // @[topLevel.scala 103:14]
  assign io_finished = co_io_finished & _T_14; // @[topLevel.scala 90:15]
  assign cfm_clock = clock;
  assign cfm_reset = reset;
  assign cfm_io_start = io_start & _T; // @[topLevel.scala 83:16]
  assign cfm_io_input_dataIn_0 = io_characterFrequencyInputs_dataIn_0; // @[topLevel.scala 93:31]
  assign cfm_io_input_valid = io_characterFrequencyInputs_valid; // @[topLevel.scala 93:31]
  assign tg_clock = clock;
  assign tg_reset = reset;
  assign tg_io_start = cfm_io_finished & _T_2; // @[topLevel.scala 84:15]
  assign tg_io_inputs_sortedFrequency_0 = cfm_io_outputs_sortedFrequency_0; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_1 = cfm_io_outputs_sortedFrequency_1; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_2 = cfm_io_outputs_sortedFrequency_2; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_3 = cfm_io_outputs_sortedFrequency_3; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_4 = cfm_io_outputs_sortedFrequency_4; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_5 = cfm_io_outputs_sortedFrequency_5; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_6 = cfm_io_outputs_sortedFrequency_6; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_7 = cfm_io_outputs_sortedFrequency_7; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_8 = cfm_io_outputs_sortedFrequency_8; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_9 = cfm_io_outputs_sortedFrequency_9; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_10 = cfm_io_outputs_sortedFrequency_10; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_11 = cfm_io_outputs_sortedFrequency_11; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_12 = cfm_io_outputs_sortedFrequency_12; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_13 = cfm_io_outputs_sortedFrequency_13; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_14 = cfm_io_outputs_sortedFrequency_14; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_15 = cfm_io_outputs_sortedFrequency_15; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_16 = cfm_io_outputs_sortedFrequency_16; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_17 = cfm_io_outputs_sortedFrequency_17; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_18 = cfm_io_outputs_sortedFrequency_18; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_19 = cfm_io_outputs_sortedFrequency_19; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_20 = cfm_io_outputs_sortedFrequency_20; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_21 = cfm_io_outputs_sortedFrequency_21; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_22 = cfm_io_outputs_sortedFrequency_22; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_23 = cfm_io_outputs_sortedFrequency_23; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_24 = cfm_io_outputs_sortedFrequency_24; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_25 = cfm_io_outputs_sortedFrequency_25; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_26 = cfm_io_outputs_sortedFrequency_26; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_27 = cfm_io_outputs_sortedFrequency_27; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_28 = cfm_io_outputs_sortedFrequency_28; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_29 = cfm_io_outputs_sortedFrequency_29; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_30 = cfm_io_outputs_sortedFrequency_30; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedFrequency_31 = cfm_io_outputs_sortedFrequency_31; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_0 = cfm_io_outputs_sortedCharacter_0; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_1 = cfm_io_outputs_sortedCharacter_1; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_2 = cfm_io_outputs_sortedCharacter_2; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_3 = cfm_io_outputs_sortedCharacter_3; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_4 = cfm_io_outputs_sortedCharacter_4; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_5 = cfm_io_outputs_sortedCharacter_5; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_6 = cfm_io_outputs_sortedCharacter_6; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_7 = cfm_io_outputs_sortedCharacter_7; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_8 = cfm_io_outputs_sortedCharacter_8; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_9 = cfm_io_outputs_sortedCharacter_9; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_10 = cfm_io_outputs_sortedCharacter_10; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_11 = cfm_io_outputs_sortedCharacter_11; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_12 = cfm_io_outputs_sortedCharacter_12; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_13 = cfm_io_outputs_sortedCharacter_13; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_14 = cfm_io_outputs_sortedCharacter_14; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_15 = cfm_io_outputs_sortedCharacter_15; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_16 = cfm_io_outputs_sortedCharacter_16; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_17 = cfm_io_outputs_sortedCharacter_17; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_18 = cfm_io_outputs_sortedCharacter_18; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_19 = cfm_io_outputs_sortedCharacter_19; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_20 = cfm_io_outputs_sortedCharacter_20; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_21 = cfm_io_outputs_sortedCharacter_21; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_22 = cfm_io_outputs_sortedCharacter_22; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_23 = cfm_io_outputs_sortedCharacter_23; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_24 = cfm_io_outputs_sortedCharacter_24; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_25 = cfm_io_outputs_sortedCharacter_25; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_26 = cfm_io_outputs_sortedCharacter_26; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_27 = cfm_io_outputs_sortedCharacter_27; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_28 = cfm_io_outputs_sortedCharacter_28; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_29 = cfm_io_outputs_sortedCharacter_29; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_30 = cfm_io_outputs_sortedCharacter_30; // @[topLevel.scala 97:16]
  assign tg_io_inputs_sortedCharacter_31 = cfm_io_outputs_sortedCharacter_31; // @[topLevel.scala 97:16]
  assign tdc_clock = clock;
  assign tdc_reset = reset;
  assign tdc_io_start = tg_io_finished & _T_4; // @[topLevel.scala 85:16]
  assign tdc_io_inputs_leftNode_0 = tg_io_outputs_leftNode_0; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_1 = tg_io_outputs_leftNode_1; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_2 = tg_io_outputs_leftNode_2; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_3 = tg_io_outputs_leftNode_3; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_4 = tg_io_outputs_leftNode_4; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_5 = tg_io_outputs_leftNode_5; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_6 = tg_io_outputs_leftNode_6; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_7 = tg_io_outputs_leftNode_7; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_8 = tg_io_outputs_leftNode_8; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_9 = tg_io_outputs_leftNode_9; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_10 = tg_io_outputs_leftNode_10; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_11 = tg_io_outputs_leftNode_11; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_12 = tg_io_outputs_leftNode_12; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_13 = tg_io_outputs_leftNode_13; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_14 = tg_io_outputs_leftNode_14; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_15 = tg_io_outputs_leftNode_15; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_16 = tg_io_outputs_leftNode_16; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_17 = tg_io_outputs_leftNode_17; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_18 = tg_io_outputs_leftNode_18; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_19 = tg_io_outputs_leftNode_19; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_20 = tg_io_outputs_leftNode_20; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_21 = tg_io_outputs_leftNode_21; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_22 = tg_io_outputs_leftNode_22; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_23 = tg_io_outputs_leftNode_23; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_24 = tg_io_outputs_leftNode_24; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_25 = tg_io_outputs_leftNode_25; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_26 = tg_io_outputs_leftNode_26; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_27 = tg_io_outputs_leftNode_27; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_28 = tg_io_outputs_leftNode_28; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_29 = tg_io_outputs_leftNode_29; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_30 = tg_io_outputs_leftNode_30; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_31 = tg_io_outputs_leftNode_31; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_32 = tg_io_outputs_leftNode_32; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_33 = tg_io_outputs_leftNode_33; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_34 = tg_io_outputs_leftNode_34; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_35 = tg_io_outputs_leftNode_35; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_36 = tg_io_outputs_leftNode_36; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_37 = tg_io_outputs_leftNode_37; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_38 = tg_io_outputs_leftNode_38; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_39 = tg_io_outputs_leftNode_39; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_40 = tg_io_outputs_leftNode_40; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_41 = tg_io_outputs_leftNode_41; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_42 = tg_io_outputs_leftNode_42; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_43 = tg_io_outputs_leftNode_43; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_44 = tg_io_outputs_leftNode_44; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_45 = tg_io_outputs_leftNode_45; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_46 = tg_io_outputs_leftNode_46; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_47 = tg_io_outputs_leftNode_47; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_48 = tg_io_outputs_leftNode_48; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_49 = tg_io_outputs_leftNode_49; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_50 = tg_io_outputs_leftNode_50; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_51 = tg_io_outputs_leftNode_51; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_52 = tg_io_outputs_leftNode_52; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_53 = tg_io_outputs_leftNode_53; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_54 = tg_io_outputs_leftNode_54; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_55 = tg_io_outputs_leftNode_55; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_56 = tg_io_outputs_leftNode_56; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_57 = tg_io_outputs_leftNode_57; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_58 = tg_io_outputs_leftNode_58; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_59 = tg_io_outputs_leftNode_59; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_60 = tg_io_outputs_leftNode_60; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_61 = tg_io_outputs_leftNode_61; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_62 = tg_io_outputs_leftNode_62; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNode_63 = tg_io_outputs_leftNode_63; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_0 = tg_io_outputs_rightNode_0; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_1 = tg_io_outputs_rightNode_1; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_2 = tg_io_outputs_rightNode_2; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_3 = tg_io_outputs_rightNode_3; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_4 = tg_io_outputs_rightNode_4; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_5 = tg_io_outputs_rightNode_5; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_6 = tg_io_outputs_rightNode_6; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_7 = tg_io_outputs_rightNode_7; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_8 = tg_io_outputs_rightNode_8; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_9 = tg_io_outputs_rightNode_9; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_10 = tg_io_outputs_rightNode_10; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_11 = tg_io_outputs_rightNode_11; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_12 = tg_io_outputs_rightNode_12; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_13 = tg_io_outputs_rightNode_13; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_14 = tg_io_outputs_rightNode_14; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_15 = tg_io_outputs_rightNode_15; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_16 = tg_io_outputs_rightNode_16; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_17 = tg_io_outputs_rightNode_17; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_18 = tg_io_outputs_rightNode_18; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_19 = tg_io_outputs_rightNode_19; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_20 = tg_io_outputs_rightNode_20; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_21 = tg_io_outputs_rightNode_21; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_22 = tg_io_outputs_rightNode_22; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_23 = tg_io_outputs_rightNode_23; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_24 = tg_io_outputs_rightNode_24; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_25 = tg_io_outputs_rightNode_25; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_26 = tg_io_outputs_rightNode_26; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_27 = tg_io_outputs_rightNode_27; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_28 = tg_io_outputs_rightNode_28; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_29 = tg_io_outputs_rightNode_29; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_30 = tg_io_outputs_rightNode_30; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_31 = tg_io_outputs_rightNode_31; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_32 = tg_io_outputs_rightNode_32; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_33 = tg_io_outputs_rightNode_33; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_34 = tg_io_outputs_rightNode_34; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_35 = tg_io_outputs_rightNode_35; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_36 = tg_io_outputs_rightNode_36; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_37 = tg_io_outputs_rightNode_37; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_38 = tg_io_outputs_rightNode_38; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_39 = tg_io_outputs_rightNode_39; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_40 = tg_io_outputs_rightNode_40; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_41 = tg_io_outputs_rightNode_41; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_42 = tg_io_outputs_rightNode_42; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_43 = tg_io_outputs_rightNode_43; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_44 = tg_io_outputs_rightNode_44; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_45 = tg_io_outputs_rightNode_45; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_46 = tg_io_outputs_rightNode_46; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_47 = tg_io_outputs_rightNode_47; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_48 = tg_io_outputs_rightNode_48; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_49 = tg_io_outputs_rightNode_49; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_50 = tg_io_outputs_rightNode_50; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_51 = tg_io_outputs_rightNode_51; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_52 = tg_io_outputs_rightNode_52; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_53 = tg_io_outputs_rightNode_53; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_54 = tg_io_outputs_rightNode_54; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_55 = tg_io_outputs_rightNode_55; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_56 = tg_io_outputs_rightNode_56; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_57 = tg_io_outputs_rightNode_57; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_58 = tg_io_outputs_rightNode_58; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_59 = tg_io_outputs_rightNode_59; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_60 = tg_io_outputs_rightNode_60; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_61 = tg_io_outputs_rightNode_61; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_62 = tg_io_outputs_rightNode_62; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNode_63 = tg_io_outputs_rightNode_63; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_0 = tg_io_outputs_leftNodeIsCharacter_0; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_1 = tg_io_outputs_leftNodeIsCharacter_1; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_2 = tg_io_outputs_leftNodeIsCharacter_2; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_3 = tg_io_outputs_leftNodeIsCharacter_3; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_4 = tg_io_outputs_leftNodeIsCharacter_4; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_5 = tg_io_outputs_leftNodeIsCharacter_5; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_6 = tg_io_outputs_leftNodeIsCharacter_6; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_7 = tg_io_outputs_leftNodeIsCharacter_7; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_8 = tg_io_outputs_leftNodeIsCharacter_8; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_9 = tg_io_outputs_leftNodeIsCharacter_9; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_10 = tg_io_outputs_leftNodeIsCharacter_10; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_11 = tg_io_outputs_leftNodeIsCharacter_11; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_12 = tg_io_outputs_leftNodeIsCharacter_12; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_13 = tg_io_outputs_leftNodeIsCharacter_13; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_14 = tg_io_outputs_leftNodeIsCharacter_14; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_15 = tg_io_outputs_leftNodeIsCharacter_15; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_16 = tg_io_outputs_leftNodeIsCharacter_16; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_17 = tg_io_outputs_leftNodeIsCharacter_17; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_18 = tg_io_outputs_leftNodeIsCharacter_18; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_19 = tg_io_outputs_leftNodeIsCharacter_19; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_20 = tg_io_outputs_leftNodeIsCharacter_20; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_21 = tg_io_outputs_leftNodeIsCharacter_21; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_22 = tg_io_outputs_leftNodeIsCharacter_22; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_23 = tg_io_outputs_leftNodeIsCharacter_23; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_24 = tg_io_outputs_leftNodeIsCharacter_24; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_25 = tg_io_outputs_leftNodeIsCharacter_25; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_26 = tg_io_outputs_leftNodeIsCharacter_26; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_27 = tg_io_outputs_leftNodeIsCharacter_27; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_28 = tg_io_outputs_leftNodeIsCharacter_28; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_29 = tg_io_outputs_leftNodeIsCharacter_29; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_30 = tg_io_outputs_leftNodeIsCharacter_30; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_31 = tg_io_outputs_leftNodeIsCharacter_31; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_32 = tg_io_outputs_leftNodeIsCharacter_32; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_33 = tg_io_outputs_leftNodeIsCharacter_33; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_34 = tg_io_outputs_leftNodeIsCharacter_34; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_35 = tg_io_outputs_leftNodeIsCharacter_35; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_36 = tg_io_outputs_leftNodeIsCharacter_36; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_37 = tg_io_outputs_leftNodeIsCharacter_37; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_38 = tg_io_outputs_leftNodeIsCharacter_38; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_39 = tg_io_outputs_leftNodeIsCharacter_39; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_40 = tg_io_outputs_leftNodeIsCharacter_40; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_41 = tg_io_outputs_leftNodeIsCharacter_41; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_42 = tg_io_outputs_leftNodeIsCharacter_42; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_43 = tg_io_outputs_leftNodeIsCharacter_43; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_44 = tg_io_outputs_leftNodeIsCharacter_44; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_45 = tg_io_outputs_leftNodeIsCharacter_45; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_46 = tg_io_outputs_leftNodeIsCharacter_46; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_47 = tg_io_outputs_leftNodeIsCharacter_47; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_48 = tg_io_outputs_leftNodeIsCharacter_48; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_49 = tg_io_outputs_leftNodeIsCharacter_49; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_50 = tg_io_outputs_leftNodeIsCharacter_50; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_51 = tg_io_outputs_leftNodeIsCharacter_51; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_52 = tg_io_outputs_leftNodeIsCharacter_52; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_53 = tg_io_outputs_leftNodeIsCharacter_53; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_54 = tg_io_outputs_leftNodeIsCharacter_54; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_55 = tg_io_outputs_leftNodeIsCharacter_55; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_56 = tg_io_outputs_leftNodeIsCharacter_56; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_57 = tg_io_outputs_leftNodeIsCharacter_57; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_58 = tg_io_outputs_leftNodeIsCharacter_58; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_59 = tg_io_outputs_leftNodeIsCharacter_59; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_60 = tg_io_outputs_leftNodeIsCharacter_60; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_61 = tg_io_outputs_leftNodeIsCharacter_61; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_62 = tg_io_outputs_leftNodeIsCharacter_62; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_leftNodeIsCharacter_63 = tg_io_outputs_leftNodeIsCharacter_63; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_0 = tg_io_outputs_rightNodeIsCharacter_0; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_1 = tg_io_outputs_rightNodeIsCharacter_1; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_2 = tg_io_outputs_rightNodeIsCharacter_2; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_3 = tg_io_outputs_rightNodeIsCharacter_3; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_4 = tg_io_outputs_rightNodeIsCharacter_4; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_5 = tg_io_outputs_rightNodeIsCharacter_5; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_6 = tg_io_outputs_rightNodeIsCharacter_6; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_7 = tg_io_outputs_rightNodeIsCharacter_7; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_8 = tg_io_outputs_rightNodeIsCharacter_8; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_9 = tg_io_outputs_rightNodeIsCharacter_9; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_10 = tg_io_outputs_rightNodeIsCharacter_10; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_11 = tg_io_outputs_rightNodeIsCharacter_11; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_12 = tg_io_outputs_rightNodeIsCharacter_12; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_13 = tg_io_outputs_rightNodeIsCharacter_13; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_14 = tg_io_outputs_rightNodeIsCharacter_14; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_15 = tg_io_outputs_rightNodeIsCharacter_15; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_16 = tg_io_outputs_rightNodeIsCharacter_16; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_17 = tg_io_outputs_rightNodeIsCharacter_17; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_18 = tg_io_outputs_rightNodeIsCharacter_18; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_19 = tg_io_outputs_rightNodeIsCharacter_19; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_20 = tg_io_outputs_rightNodeIsCharacter_20; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_21 = tg_io_outputs_rightNodeIsCharacter_21; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_22 = tg_io_outputs_rightNodeIsCharacter_22; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_23 = tg_io_outputs_rightNodeIsCharacter_23; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_24 = tg_io_outputs_rightNodeIsCharacter_24; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_25 = tg_io_outputs_rightNodeIsCharacter_25; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_26 = tg_io_outputs_rightNodeIsCharacter_26; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_27 = tg_io_outputs_rightNodeIsCharacter_27; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_28 = tg_io_outputs_rightNodeIsCharacter_28; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_29 = tg_io_outputs_rightNodeIsCharacter_29; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_30 = tg_io_outputs_rightNodeIsCharacter_30; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_31 = tg_io_outputs_rightNodeIsCharacter_31; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_32 = tg_io_outputs_rightNodeIsCharacter_32; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_33 = tg_io_outputs_rightNodeIsCharacter_33; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_34 = tg_io_outputs_rightNodeIsCharacter_34; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_35 = tg_io_outputs_rightNodeIsCharacter_35; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_36 = tg_io_outputs_rightNodeIsCharacter_36; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_37 = tg_io_outputs_rightNodeIsCharacter_37; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_38 = tg_io_outputs_rightNodeIsCharacter_38; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_39 = tg_io_outputs_rightNodeIsCharacter_39; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_40 = tg_io_outputs_rightNodeIsCharacter_40; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_41 = tg_io_outputs_rightNodeIsCharacter_41; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_42 = tg_io_outputs_rightNodeIsCharacter_42; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_43 = tg_io_outputs_rightNodeIsCharacter_43; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_44 = tg_io_outputs_rightNodeIsCharacter_44; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_45 = tg_io_outputs_rightNodeIsCharacter_45; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_46 = tg_io_outputs_rightNodeIsCharacter_46; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_47 = tg_io_outputs_rightNodeIsCharacter_47; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_48 = tg_io_outputs_rightNodeIsCharacter_48; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_49 = tg_io_outputs_rightNodeIsCharacter_49; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_50 = tg_io_outputs_rightNodeIsCharacter_50; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_51 = tg_io_outputs_rightNodeIsCharacter_51; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_52 = tg_io_outputs_rightNodeIsCharacter_52; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_53 = tg_io_outputs_rightNodeIsCharacter_53; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_54 = tg_io_outputs_rightNodeIsCharacter_54; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_55 = tg_io_outputs_rightNodeIsCharacter_55; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_56 = tg_io_outputs_rightNodeIsCharacter_56; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_57 = tg_io_outputs_rightNodeIsCharacter_57; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_58 = tg_io_outputs_rightNodeIsCharacter_58; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_59 = tg_io_outputs_rightNodeIsCharacter_59; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_60 = tg_io_outputs_rightNodeIsCharacter_60; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_61 = tg_io_outputs_rightNodeIsCharacter_61; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_62 = tg_io_outputs_rightNodeIsCharacter_62; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_rightNodeIsCharacter_63 = tg_io_outputs_rightNodeIsCharacter_63; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_validNodes = tg_io_outputs_validNodes; // @[topLevel.scala 98:17]
  assign tdc_io_inputs_validCharacters = tg_io_outputs_validCharacters; // @[topLevel.scala 98:17]
  assign sltg_clock = clock;
  assign sltg_reset = reset;
  assign sltg_io_start = tdc_io_finished & _T_6; // @[topLevel.scala 86:17]
  assign sltg_io_inputs_characters_0 = tdc_io_outputs_characters_0; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_1 = tdc_io_outputs_characters_1; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_2 = tdc_io_outputs_characters_2; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_3 = tdc_io_outputs_characters_3; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_4 = tdc_io_outputs_characters_4; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_5 = tdc_io_outputs_characters_5; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_6 = tdc_io_outputs_characters_6; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_7 = tdc_io_outputs_characters_7; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_8 = tdc_io_outputs_characters_8; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_9 = tdc_io_outputs_characters_9; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_10 = tdc_io_outputs_characters_10; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_11 = tdc_io_outputs_characters_11; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_12 = tdc_io_outputs_characters_12; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_13 = tdc_io_outputs_characters_13; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_14 = tdc_io_outputs_characters_14; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_15 = tdc_io_outputs_characters_15; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_16 = tdc_io_outputs_characters_16; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_17 = tdc_io_outputs_characters_17; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_18 = tdc_io_outputs_characters_18; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_19 = tdc_io_outputs_characters_19; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_20 = tdc_io_outputs_characters_20; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_21 = tdc_io_outputs_characters_21; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_22 = tdc_io_outputs_characters_22; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_23 = tdc_io_outputs_characters_23; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_24 = tdc_io_outputs_characters_24; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_25 = tdc_io_outputs_characters_25; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_26 = tdc_io_outputs_characters_26; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_27 = tdc_io_outputs_characters_27; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_28 = tdc_io_outputs_characters_28; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_29 = tdc_io_outputs_characters_29; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_30 = tdc_io_outputs_characters_30; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_characters_31 = tdc_io_outputs_characters_31; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_0 = tdc_io_outputs_depths_0; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_1 = tdc_io_outputs_depths_1; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_2 = tdc_io_outputs_depths_2; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_3 = tdc_io_outputs_depths_3; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_4 = tdc_io_outputs_depths_4; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_5 = tdc_io_outputs_depths_5; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_6 = tdc_io_outputs_depths_6; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_7 = tdc_io_outputs_depths_7; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_8 = tdc_io_outputs_depths_8; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_9 = tdc_io_outputs_depths_9; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_10 = tdc_io_outputs_depths_10; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_11 = tdc_io_outputs_depths_11; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_12 = tdc_io_outputs_depths_12; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_13 = tdc_io_outputs_depths_13; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_14 = tdc_io_outputs_depths_14; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_15 = tdc_io_outputs_depths_15; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_16 = tdc_io_outputs_depths_16; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_17 = tdc_io_outputs_depths_17; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_18 = tdc_io_outputs_depths_18; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_19 = tdc_io_outputs_depths_19; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_20 = tdc_io_outputs_depths_20; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_21 = tdc_io_outputs_depths_21; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_22 = tdc_io_outputs_depths_22; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_23 = tdc_io_outputs_depths_23; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_24 = tdc_io_outputs_depths_24; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_25 = tdc_io_outputs_depths_25; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_26 = tdc_io_outputs_depths_26; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_27 = tdc_io_outputs_depths_27; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_28 = tdc_io_outputs_depths_28; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_29 = tdc_io_outputs_depths_29; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_30 = tdc_io_outputs_depths_30; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_depths_31 = tdc_io_outputs_depths_31; // @[topLevel.scala 99:18]
  assign sltg_io_inputs_validCharacters = tdc_io_outputs_validCharacters; // @[topLevel.scala 99:18]
  assign tn_clock = clock;
  assign tn_reset = reset;
  assign tn_io_start = sltg_io_finished & _T_8; // @[topLevel.scala 87:15]
  assign tn_io_inputs_outputData_0 = sltg_io_outputs_outputData_0; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_1 = sltg_io_outputs_outputData_1; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_2 = sltg_io_outputs_outputData_2; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_3 = sltg_io_outputs_outputData_3; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_4 = sltg_io_outputs_outputData_4; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_5 = sltg_io_outputs_outputData_5; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_6 = sltg_io_outputs_outputData_6; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_7 = sltg_io_outputs_outputData_7; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_8 = sltg_io_outputs_outputData_8; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_9 = sltg_io_outputs_outputData_9; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_10 = sltg_io_outputs_outputData_10; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_11 = sltg_io_outputs_outputData_11; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_12 = sltg_io_outputs_outputData_12; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_13 = sltg_io_outputs_outputData_13; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_14 = sltg_io_outputs_outputData_14; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_15 = sltg_io_outputs_outputData_15; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_16 = sltg_io_outputs_outputData_16; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_17 = sltg_io_outputs_outputData_17; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_18 = sltg_io_outputs_outputData_18; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_19 = sltg_io_outputs_outputData_19; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_20 = sltg_io_outputs_outputData_20; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_21 = sltg_io_outputs_outputData_21; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_22 = sltg_io_outputs_outputData_22; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_23 = sltg_io_outputs_outputData_23; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_24 = sltg_io_outputs_outputData_24; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_25 = sltg_io_outputs_outputData_25; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_26 = sltg_io_outputs_outputData_26; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_27 = sltg_io_outputs_outputData_27; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_28 = sltg_io_outputs_outputData_28; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_29 = sltg_io_outputs_outputData_29; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_30 = sltg_io_outputs_outputData_30; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputData_31 = sltg_io_outputs_outputData_31; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_0 = sltg_io_outputs_outputTags_0; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_1 = sltg_io_outputs_outputTags_1; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_2 = sltg_io_outputs_outputTags_2; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_3 = sltg_io_outputs_outputTags_3; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_4 = sltg_io_outputs_outputTags_4; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_5 = sltg_io_outputs_outputTags_5; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_6 = sltg_io_outputs_outputTags_6; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_7 = sltg_io_outputs_outputTags_7; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_8 = sltg_io_outputs_outputTags_8; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_9 = sltg_io_outputs_outputTags_9; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_10 = sltg_io_outputs_outputTags_10; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_11 = sltg_io_outputs_outputTags_11; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_12 = sltg_io_outputs_outputTags_12; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_13 = sltg_io_outputs_outputTags_13; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_14 = sltg_io_outputs_outputTags_14; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_15 = sltg_io_outputs_outputTags_15; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_16 = sltg_io_outputs_outputTags_16; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_17 = sltg_io_outputs_outputTags_17; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_18 = sltg_io_outputs_outputTags_18; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_19 = sltg_io_outputs_outputTags_19; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_20 = sltg_io_outputs_outputTags_20; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_21 = sltg_io_outputs_outputTags_21; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_22 = sltg_io_outputs_outputTags_22; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_23 = sltg_io_outputs_outputTags_23; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_24 = sltg_io_outputs_outputTags_24; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_25 = sltg_io_outputs_outputTags_25; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_26 = sltg_io_outputs_outputTags_26; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_27 = sltg_io_outputs_outputTags_27; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_28 = sltg_io_outputs_outputTags_28; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_29 = sltg_io_outputs_outputTags_29; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_30 = sltg_io_outputs_outputTags_30; // @[topLevel.scala 100:16]
  assign tn_io_inputs_outputTags_31 = sltg_io_outputs_outputTags_31; // @[topLevel.scala 100:16]
  assign tn_io_inputs_itemNumber = sltg_io_outputs_itemNumber; // @[topLevel.scala 100:16]
  assign cg_clock = clock;
  assign cg_reset = reset;
  assign cg_io_start = tn_io_finished & _T_10; // @[topLevel.scala 88:15]
  assign cg_io_inputs_charactersOut_0 = tn_io_outputs_charactersOut_0; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_1 = tn_io_outputs_charactersOut_1; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_2 = tn_io_outputs_charactersOut_2; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_3 = tn_io_outputs_charactersOut_3; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_4 = tn_io_outputs_charactersOut_4; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_5 = tn_io_outputs_charactersOut_5; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_6 = tn_io_outputs_charactersOut_6; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_7 = tn_io_outputs_charactersOut_7; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_8 = tn_io_outputs_charactersOut_8; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_9 = tn_io_outputs_charactersOut_9; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_10 = tn_io_outputs_charactersOut_10; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_11 = tn_io_outputs_charactersOut_11; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_12 = tn_io_outputs_charactersOut_12; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_13 = tn_io_outputs_charactersOut_13; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_14 = tn_io_outputs_charactersOut_14; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_15 = tn_io_outputs_charactersOut_15; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_16 = tn_io_outputs_charactersOut_16; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_17 = tn_io_outputs_charactersOut_17; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_18 = tn_io_outputs_charactersOut_18; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_19 = tn_io_outputs_charactersOut_19; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_20 = tn_io_outputs_charactersOut_20; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_21 = tn_io_outputs_charactersOut_21; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_22 = tn_io_outputs_charactersOut_22; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_23 = tn_io_outputs_charactersOut_23; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_24 = tn_io_outputs_charactersOut_24; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_25 = tn_io_outputs_charactersOut_25; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_26 = tn_io_outputs_charactersOut_26; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_27 = tn_io_outputs_charactersOut_27; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_28 = tn_io_outputs_charactersOut_28; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_29 = tn_io_outputs_charactersOut_29; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_30 = tn_io_outputs_charactersOut_30; // @[topLevel.scala 101:16]
  assign cg_io_inputs_charactersOut_31 = tn_io_outputs_charactersOut_31; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_0 = tn_io_outputs_depthsOut_0; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_1 = tn_io_outputs_depthsOut_1; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_2 = tn_io_outputs_depthsOut_2; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_3 = tn_io_outputs_depthsOut_3; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_4 = tn_io_outputs_depthsOut_4; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_5 = tn_io_outputs_depthsOut_5; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_6 = tn_io_outputs_depthsOut_6; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_7 = tn_io_outputs_depthsOut_7; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_8 = tn_io_outputs_depthsOut_8; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_9 = tn_io_outputs_depthsOut_9; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_10 = tn_io_outputs_depthsOut_10; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_11 = tn_io_outputs_depthsOut_11; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_12 = tn_io_outputs_depthsOut_12; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_13 = tn_io_outputs_depthsOut_13; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_14 = tn_io_outputs_depthsOut_14; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_15 = tn_io_outputs_depthsOut_15; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_16 = tn_io_outputs_depthsOut_16; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_17 = tn_io_outputs_depthsOut_17; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_18 = tn_io_outputs_depthsOut_18; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_19 = tn_io_outputs_depthsOut_19; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_20 = tn_io_outputs_depthsOut_20; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_21 = tn_io_outputs_depthsOut_21; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_22 = tn_io_outputs_depthsOut_22; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_23 = tn_io_outputs_depthsOut_23; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_24 = tn_io_outputs_depthsOut_24; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_25 = tn_io_outputs_depthsOut_25; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_26 = tn_io_outputs_depthsOut_26; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_27 = tn_io_outputs_depthsOut_27; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_28 = tn_io_outputs_depthsOut_28; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_29 = tn_io_outputs_depthsOut_29; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_30 = tn_io_outputs_depthsOut_30; // @[topLevel.scala 101:16]
  assign cg_io_inputs_depthsOut_31 = tn_io_outputs_depthsOut_31; // @[topLevel.scala 101:16]
  assign cg_io_inputs_validNodesOut = tn_io_outputs_validNodesOut; // @[topLevel.scala 101:16]
  assign co_clock = clock;
  assign co_reset = reset;
  assign co_io_start = cg_io_finished & _T_12; // @[topLevel.scala 89:15]
  assign co_io_dataIn_0_dataIn_0 = io_compressionInputs_0_dataIn_0; // @[topLevel.scala 95:33]
  assign co_io_dataIn_0_valid = io_compressionInputs_0_valid; // @[topLevel.scala 95:33]
  assign co_io_inputs_codewords_0 = cg_io_outputs_codewords_0; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_1 = cg_io_outputs_codewords_1; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_2 = cg_io_outputs_codewords_2; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_3 = cg_io_outputs_codewords_3; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_4 = cg_io_outputs_codewords_4; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_5 = cg_io_outputs_codewords_5; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_6 = cg_io_outputs_codewords_6; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_7 = cg_io_outputs_codewords_7; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_8 = cg_io_outputs_codewords_8; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_9 = cg_io_outputs_codewords_9; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_10 = cg_io_outputs_codewords_10; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_11 = cg_io_outputs_codewords_11; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_12 = cg_io_outputs_codewords_12; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_13 = cg_io_outputs_codewords_13; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_14 = cg_io_outputs_codewords_14; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_15 = cg_io_outputs_codewords_15; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_16 = cg_io_outputs_codewords_16; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_17 = cg_io_outputs_codewords_17; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_18 = cg_io_outputs_codewords_18; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_19 = cg_io_outputs_codewords_19; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_20 = cg_io_outputs_codewords_20; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_21 = cg_io_outputs_codewords_21; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_22 = cg_io_outputs_codewords_22; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_23 = cg_io_outputs_codewords_23; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_24 = cg_io_outputs_codewords_24; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_25 = cg_io_outputs_codewords_25; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_26 = cg_io_outputs_codewords_26; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_27 = cg_io_outputs_codewords_27; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_28 = cg_io_outputs_codewords_28; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_29 = cg_io_outputs_codewords_29; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_30 = cg_io_outputs_codewords_30; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_31 = cg_io_outputs_codewords_31; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_32 = cg_io_outputs_codewords_32; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_33 = cg_io_outputs_codewords_33; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_34 = cg_io_outputs_codewords_34; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_35 = cg_io_outputs_codewords_35; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_36 = cg_io_outputs_codewords_36; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_37 = cg_io_outputs_codewords_37; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_38 = cg_io_outputs_codewords_38; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_39 = cg_io_outputs_codewords_39; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_40 = cg_io_outputs_codewords_40; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_41 = cg_io_outputs_codewords_41; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_42 = cg_io_outputs_codewords_42; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_43 = cg_io_outputs_codewords_43; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_44 = cg_io_outputs_codewords_44; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_45 = cg_io_outputs_codewords_45; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_46 = cg_io_outputs_codewords_46; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_47 = cg_io_outputs_codewords_47; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_48 = cg_io_outputs_codewords_48; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_49 = cg_io_outputs_codewords_49; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_50 = cg_io_outputs_codewords_50; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_51 = cg_io_outputs_codewords_51; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_52 = cg_io_outputs_codewords_52; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_53 = cg_io_outputs_codewords_53; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_54 = cg_io_outputs_codewords_54; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_55 = cg_io_outputs_codewords_55; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_56 = cg_io_outputs_codewords_56; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_57 = cg_io_outputs_codewords_57; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_58 = cg_io_outputs_codewords_58; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_59 = cg_io_outputs_codewords_59; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_60 = cg_io_outputs_codewords_60; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_61 = cg_io_outputs_codewords_61; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_62 = cg_io_outputs_codewords_62; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_63 = cg_io_outputs_codewords_63; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_64 = cg_io_outputs_codewords_64; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_65 = cg_io_outputs_codewords_65; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_66 = cg_io_outputs_codewords_66; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_67 = cg_io_outputs_codewords_67; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_68 = cg_io_outputs_codewords_68; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_69 = cg_io_outputs_codewords_69; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_70 = cg_io_outputs_codewords_70; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_71 = cg_io_outputs_codewords_71; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_72 = cg_io_outputs_codewords_72; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_73 = cg_io_outputs_codewords_73; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_74 = cg_io_outputs_codewords_74; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_75 = cg_io_outputs_codewords_75; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_76 = cg_io_outputs_codewords_76; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_77 = cg_io_outputs_codewords_77; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_78 = cg_io_outputs_codewords_78; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_79 = cg_io_outputs_codewords_79; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_80 = cg_io_outputs_codewords_80; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_81 = cg_io_outputs_codewords_81; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_82 = cg_io_outputs_codewords_82; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_83 = cg_io_outputs_codewords_83; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_84 = cg_io_outputs_codewords_84; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_85 = cg_io_outputs_codewords_85; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_86 = cg_io_outputs_codewords_86; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_87 = cg_io_outputs_codewords_87; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_88 = cg_io_outputs_codewords_88; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_89 = cg_io_outputs_codewords_89; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_90 = cg_io_outputs_codewords_90; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_91 = cg_io_outputs_codewords_91; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_92 = cg_io_outputs_codewords_92; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_93 = cg_io_outputs_codewords_93; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_94 = cg_io_outputs_codewords_94; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_95 = cg_io_outputs_codewords_95; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_96 = cg_io_outputs_codewords_96; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_97 = cg_io_outputs_codewords_97; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_98 = cg_io_outputs_codewords_98; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_99 = cg_io_outputs_codewords_99; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_100 = cg_io_outputs_codewords_100; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_101 = cg_io_outputs_codewords_101; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_102 = cg_io_outputs_codewords_102; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_103 = cg_io_outputs_codewords_103; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_104 = cg_io_outputs_codewords_104; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_105 = cg_io_outputs_codewords_105; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_106 = cg_io_outputs_codewords_106; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_107 = cg_io_outputs_codewords_107; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_108 = cg_io_outputs_codewords_108; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_109 = cg_io_outputs_codewords_109; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_110 = cg_io_outputs_codewords_110; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_111 = cg_io_outputs_codewords_111; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_112 = cg_io_outputs_codewords_112; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_113 = cg_io_outputs_codewords_113; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_114 = cg_io_outputs_codewords_114; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_115 = cg_io_outputs_codewords_115; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_116 = cg_io_outputs_codewords_116; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_117 = cg_io_outputs_codewords_117; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_118 = cg_io_outputs_codewords_118; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_119 = cg_io_outputs_codewords_119; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_120 = cg_io_outputs_codewords_120; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_121 = cg_io_outputs_codewords_121; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_122 = cg_io_outputs_codewords_122; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_123 = cg_io_outputs_codewords_123; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_124 = cg_io_outputs_codewords_124; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_125 = cg_io_outputs_codewords_125; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_126 = cg_io_outputs_codewords_126; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_127 = cg_io_outputs_codewords_127; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_128 = cg_io_outputs_codewords_128; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_129 = cg_io_outputs_codewords_129; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_130 = cg_io_outputs_codewords_130; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_131 = cg_io_outputs_codewords_131; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_132 = cg_io_outputs_codewords_132; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_133 = cg_io_outputs_codewords_133; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_134 = cg_io_outputs_codewords_134; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_135 = cg_io_outputs_codewords_135; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_136 = cg_io_outputs_codewords_136; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_137 = cg_io_outputs_codewords_137; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_138 = cg_io_outputs_codewords_138; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_139 = cg_io_outputs_codewords_139; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_140 = cg_io_outputs_codewords_140; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_141 = cg_io_outputs_codewords_141; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_142 = cg_io_outputs_codewords_142; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_143 = cg_io_outputs_codewords_143; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_144 = cg_io_outputs_codewords_144; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_145 = cg_io_outputs_codewords_145; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_146 = cg_io_outputs_codewords_146; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_147 = cg_io_outputs_codewords_147; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_148 = cg_io_outputs_codewords_148; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_149 = cg_io_outputs_codewords_149; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_150 = cg_io_outputs_codewords_150; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_151 = cg_io_outputs_codewords_151; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_152 = cg_io_outputs_codewords_152; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_153 = cg_io_outputs_codewords_153; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_154 = cg_io_outputs_codewords_154; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_155 = cg_io_outputs_codewords_155; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_156 = cg_io_outputs_codewords_156; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_157 = cg_io_outputs_codewords_157; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_158 = cg_io_outputs_codewords_158; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_159 = cg_io_outputs_codewords_159; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_160 = cg_io_outputs_codewords_160; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_161 = cg_io_outputs_codewords_161; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_162 = cg_io_outputs_codewords_162; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_163 = cg_io_outputs_codewords_163; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_164 = cg_io_outputs_codewords_164; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_165 = cg_io_outputs_codewords_165; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_166 = cg_io_outputs_codewords_166; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_167 = cg_io_outputs_codewords_167; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_168 = cg_io_outputs_codewords_168; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_169 = cg_io_outputs_codewords_169; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_170 = cg_io_outputs_codewords_170; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_171 = cg_io_outputs_codewords_171; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_172 = cg_io_outputs_codewords_172; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_173 = cg_io_outputs_codewords_173; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_174 = cg_io_outputs_codewords_174; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_175 = cg_io_outputs_codewords_175; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_176 = cg_io_outputs_codewords_176; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_177 = cg_io_outputs_codewords_177; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_178 = cg_io_outputs_codewords_178; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_179 = cg_io_outputs_codewords_179; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_180 = cg_io_outputs_codewords_180; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_181 = cg_io_outputs_codewords_181; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_182 = cg_io_outputs_codewords_182; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_183 = cg_io_outputs_codewords_183; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_184 = cg_io_outputs_codewords_184; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_185 = cg_io_outputs_codewords_185; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_186 = cg_io_outputs_codewords_186; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_187 = cg_io_outputs_codewords_187; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_188 = cg_io_outputs_codewords_188; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_189 = cg_io_outputs_codewords_189; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_190 = cg_io_outputs_codewords_190; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_191 = cg_io_outputs_codewords_191; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_192 = cg_io_outputs_codewords_192; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_193 = cg_io_outputs_codewords_193; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_194 = cg_io_outputs_codewords_194; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_195 = cg_io_outputs_codewords_195; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_196 = cg_io_outputs_codewords_196; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_197 = cg_io_outputs_codewords_197; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_198 = cg_io_outputs_codewords_198; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_199 = cg_io_outputs_codewords_199; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_200 = cg_io_outputs_codewords_200; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_201 = cg_io_outputs_codewords_201; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_202 = cg_io_outputs_codewords_202; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_203 = cg_io_outputs_codewords_203; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_204 = cg_io_outputs_codewords_204; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_205 = cg_io_outputs_codewords_205; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_206 = cg_io_outputs_codewords_206; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_207 = cg_io_outputs_codewords_207; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_208 = cg_io_outputs_codewords_208; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_209 = cg_io_outputs_codewords_209; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_210 = cg_io_outputs_codewords_210; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_211 = cg_io_outputs_codewords_211; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_212 = cg_io_outputs_codewords_212; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_213 = cg_io_outputs_codewords_213; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_214 = cg_io_outputs_codewords_214; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_215 = cg_io_outputs_codewords_215; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_216 = cg_io_outputs_codewords_216; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_217 = cg_io_outputs_codewords_217; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_218 = cg_io_outputs_codewords_218; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_219 = cg_io_outputs_codewords_219; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_220 = cg_io_outputs_codewords_220; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_221 = cg_io_outputs_codewords_221; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_222 = cg_io_outputs_codewords_222; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_223 = cg_io_outputs_codewords_223; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_224 = cg_io_outputs_codewords_224; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_225 = cg_io_outputs_codewords_225; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_226 = cg_io_outputs_codewords_226; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_227 = cg_io_outputs_codewords_227; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_228 = cg_io_outputs_codewords_228; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_229 = cg_io_outputs_codewords_229; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_230 = cg_io_outputs_codewords_230; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_231 = cg_io_outputs_codewords_231; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_232 = cg_io_outputs_codewords_232; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_233 = cg_io_outputs_codewords_233; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_234 = cg_io_outputs_codewords_234; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_235 = cg_io_outputs_codewords_235; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_236 = cg_io_outputs_codewords_236; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_237 = cg_io_outputs_codewords_237; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_238 = cg_io_outputs_codewords_238; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_239 = cg_io_outputs_codewords_239; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_240 = cg_io_outputs_codewords_240; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_241 = cg_io_outputs_codewords_241; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_242 = cg_io_outputs_codewords_242; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_243 = cg_io_outputs_codewords_243; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_244 = cg_io_outputs_codewords_244; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_245 = cg_io_outputs_codewords_245; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_246 = cg_io_outputs_codewords_246; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_247 = cg_io_outputs_codewords_247; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_248 = cg_io_outputs_codewords_248; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_249 = cg_io_outputs_codewords_249; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_250 = cg_io_outputs_codewords_250; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_251 = cg_io_outputs_codewords_251; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_252 = cg_io_outputs_codewords_252; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_253 = cg_io_outputs_codewords_253; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_254 = cg_io_outputs_codewords_254; // @[topLevel.scala 102:16]
  assign co_io_inputs_codewords_255 = cg_io_outputs_codewords_255; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_0 = cg_io_outputs_lengths_0; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_1 = cg_io_outputs_lengths_1; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_2 = cg_io_outputs_lengths_2; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_3 = cg_io_outputs_lengths_3; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_4 = cg_io_outputs_lengths_4; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_5 = cg_io_outputs_lengths_5; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_6 = cg_io_outputs_lengths_6; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_7 = cg_io_outputs_lengths_7; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_8 = cg_io_outputs_lengths_8; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_9 = cg_io_outputs_lengths_9; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_10 = cg_io_outputs_lengths_10; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_11 = cg_io_outputs_lengths_11; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_12 = cg_io_outputs_lengths_12; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_13 = cg_io_outputs_lengths_13; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_14 = cg_io_outputs_lengths_14; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_15 = cg_io_outputs_lengths_15; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_16 = cg_io_outputs_lengths_16; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_17 = cg_io_outputs_lengths_17; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_18 = cg_io_outputs_lengths_18; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_19 = cg_io_outputs_lengths_19; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_20 = cg_io_outputs_lengths_20; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_21 = cg_io_outputs_lengths_21; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_22 = cg_io_outputs_lengths_22; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_23 = cg_io_outputs_lengths_23; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_24 = cg_io_outputs_lengths_24; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_25 = cg_io_outputs_lengths_25; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_26 = cg_io_outputs_lengths_26; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_27 = cg_io_outputs_lengths_27; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_28 = cg_io_outputs_lengths_28; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_29 = cg_io_outputs_lengths_29; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_30 = cg_io_outputs_lengths_30; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_31 = cg_io_outputs_lengths_31; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_32 = cg_io_outputs_lengths_32; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_33 = cg_io_outputs_lengths_33; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_34 = cg_io_outputs_lengths_34; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_35 = cg_io_outputs_lengths_35; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_36 = cg_io_outputs_lengths_36; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_37 = cg_io_outputs_lengths_37; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_38 = cg_io_outputs_lengths_38; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_39 = cg_io_outputs_lengths_39; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_40 = cg_io_outputs_lengths_40; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_41 = cg_io_outputs_lengths_41; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_42 = cg_io_outputs_lengths_42; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_43 = cg_io_outputs_lengths_43; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_44 = cg_io_outputs_lengths_44; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_45 = cg_io_outputs_lengths_45; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_46 = cg_io_outputs_lengths_46; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_47 = cg_io_outputs_lengths_47; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_48 = cg_io_outputs_lengths_48; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_49 = cg_io_outputs_lengths_49; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_50 = cg_io_outputs_lengths_50; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_51 = cg_io_outputs_lengths_51; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_52 = cg_io_outputs_lengths_52; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_53 = cg_io_outputs_lengths_53; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_54 = cg_io_outputs_lengths_54; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_55 = cg_io_outputs_lengths_55; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_56 = cg_io_outputs_lengths_56; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_57 = cg_io_outputs_lengths_57; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_58 = cg_io_outputs_lengths_58; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_59 = cg_io_outputs_lengths_59; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_60 = cg_io_outputs_lengths_60; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_61 = cg_io_outputs_lengths_61; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_62 = cg_io_outputs_lengths_62; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_63 = cg_io_outputs_lengths_63; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_64 = cg_io_outputs_lengths_64; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_65 = cg_io_outputs_lengths_65; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_66 = cg_io_outputs_lengths_66; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_67 = cg_io_outputs_lengths_67; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_68 = cg_io_outputs_lengths_68; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_69 = cg_io_outputs_lengths_69; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_70 = cg_io_outputs_lengths_70; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_71 = cg_io_outputs_lengths_71; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_72 = cg_io_outputs_lengths_72; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_73 = cg_io_outputs_lengths_73; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_74 = cg_io_outputs_lengths_74; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_75 = cg_io_outputs_lengths_75; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_76 = cg_io_outputs_lengths_76; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_77 = cg_io_outputs_lengths_77; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_78 = cg_io_outputs_lengths_78; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_79 = cg_io_outputs_lengths_79; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_80 = cg_io_outputs_lengths_80; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_81 = cg_io_outputs_lengths_81; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_82 = cg_io_outputs_lengths_82; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_83 = cg_io_outputs_lengths_83; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_84 = cg_io_outputs_lengths_84; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_85 = cg_io_outputs_lengths_85; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_86 = cg_io_outputs_lengths_86; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_87 = cg_io_outputs_lengths_87; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_88 = cg_io_outputs_lengths_88; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_89 = cg_io_outputs_lengths_89; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_90 = cg_io_outputs_lengths_90; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_91 = cg_io_outputs_lengths_91; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_92 = cg_io_outputs_lengths_92; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_93 = cg_io_outputs_lengths_93; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_94 = cg_io_outputs_lengths_94; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_95 = cg_io_outputs_lengths_95; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_96 = cg_io_outputs_lengths_96; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_97 = cg_io_outputs_lengths_97; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_98 = cg_io_outputs_lengths_98; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_99 = cg_io_outputs_lengths_99; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_100 = cg_io_outputs_lengths_100; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_101 = cg_io_outputs_lengths_101; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_102 = cg_io_outputs_lengths_102; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_103 = cg_io_outputs_lengths_103; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_104 = cg_io_outputs_lengths_104; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_105 = cg_io_outputs_lengths_105; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_106 = cg_io_outputs_lengths_106; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_107 = cg_io_outputs_lengths_107; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_108 = cg_io_outputs_lengths_108; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_109 = cg_io_outputs_lengths_109; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_110 = cg_io_outputs_lengths_110; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_111 = cg_io_outputs_lengths_111; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_112 = cg_io_outputs_lengths_112; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_113 = cg_io_outputs_lengths_113; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_114 = cg_io_outputs_lengths_114; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_115 = cg_io_outputs_lengths_115; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_116 = cg_io_outputs_lengths_116; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_117 = cg_io_outputs_lengths_117; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_118 = cg_io_outputs_lengths_118; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_119 = cg_io_outputs_lengths_119; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_120 = cg_io_outputs_lengths_120; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_121 = cg_io_outputs_lengths_121; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_122 = cg_io_outputs_lengths_122; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_123 = cg_io_outputs_lengths_123; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_124 = cg_io_outputs_lengths_124; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_125 = cg_io_outputs_lengths_125; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_126 = cg_io_outputs_lengths_126; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_127 = cg_io_outputs_lengths_127; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_128 = cg_io_outputs_lengths_128; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_129 = cg_io_outputs_lengths_129; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_130 = cg_io_outputs_lengths_130; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_131 = cg_io_outputs_lengths_131; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_132 = cg_io_outputs_lengths_132; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_133 = cg_io_outputs_lengths_133; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_134 = cg_io_outputs_lengths_134; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_135 = cg_io_outputs_lengths_135; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_136 = cg_io_outputs_lengths_136; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_137 = cg_io_outputs_lengths_137; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_138 = cg_io_outputs_lengths_138; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_139 = cg_io_outputs_lengths_139; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_140 = cg_io_outputs_lengths_140; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_141 = cg_io_outputs_lengths_141; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_142 = cg_io_outputs_lengths_142; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_143 = cg_io_outputs_lengths_143; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_144 = cg_io_outputs_lengths_144; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_145 = cg_io_outputs_lengths_145; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_146 = cg_io_outputs_lengths_146; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_147 = cg_io_outputs_lengths_147; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_148 = cg_io_outputs_lengths_148; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_149 = cg_io_outputs_lengths_149; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_150 = cg_io_outputs_lengths_150; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_151 = cg_io_outputs_lengths_151; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_152 = cg_io_outputs_lengths_152; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_153 = cg_io_outputs_lengths_153; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_154 = cg_io_outputs_lengths_154; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_155 = cg_io_outputs_lengths_155; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_156 = cg_io_outputs_lengths_156; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_157 = cg_io_outputs_lengths_157; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_158 = cg_io_outputs_lengths_158; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_159 = cg_io_outputs_lengths_159; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_160 = cg_io_outputs_lengths_160; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_161 = cg_io_outputs_lengths_161; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_162 = cg_io_outputs_lengths_162; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_163 = cg_io_outputs_lengths_163; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_164 = cg_io_outputs_lengths_164; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_165 = cg_io_outputs_lengths_165; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_166 = cg_io_outputs_lengths_166; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_167 = cg_io_outputs_lengths_167; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_168 = cg_io_outputs_lengths_168; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_169 = cg_io_outputs_lengths_169; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_170 = cg_io_outputs_lengths_170; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_171 = cg_io_outputs_lengths_171; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_172 = cg_io_outputs_lengths_172; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_173 = cg_io_outputs_lengths_173; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_174 = cg_io_outputs_lengths_174; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_175 = cg_io_outputs_lengths_175; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_176 = cg_io_outputs_lengths_176; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_177 = cg_io_outputs_lengths_177; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_178 = cg_io_outputs_lengths_178; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_179 = cg_io_outputs_lengths_179; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_180 = cg_io_outputs_lengths_180; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_181 = cg_io_outputs_lengths_181; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_182 = cg_io_outputs_lengths_182; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_183 = cg_io_outputs_lengths_183; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_184 = cg_io_outputs_lengths_184; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_185 = cg_io_outputs_lengths_185; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_186 = cg_io_outputs_lengths_186; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_187 = cg_io_outputs_lengths_187; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_188 = cg_io_outputs_lengths_188; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_189 = cg_io_outputs_lengths_189; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_190 = cg_io_outputs_lengths_190; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_191 = cg_io_outputs_lengths_191; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_192 = cg_io_outputs_lengths_192; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_193 = cg_io_outputs_lengths_193; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_194 = cg_io_outputs_lengths_194; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_195 = cg_io_outputs_lengths_195; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_196 = cg_io_outputs_lengths_196; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_197 = cg_io_outputs_lengths_197; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_198 = cg_io_outputs_lengths_198; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_199 = cg_io_outputs_lengths_199; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_200 = cg_io_outputs_lengths_200; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_201 = cg_io_outputs_lengths_201; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_202 = cg_io_outputs_lengths_202; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_203 = cg_io_outputs_lengths_203; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_204 = cg_io_outputs_lengths_204; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_205 = cg_io_outputs_lengths_205; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_206 = cg_io_outputs_lengths_206; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_207 = cg_io_outputs_lengths_207; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_208 = cg_io_outputs_lengths_208; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_209 = cg_io_outputs_lengths_209; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_210 = cg_io_outputs_lengths_210; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_211 = cg_io_outputs_lengths_211; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_212 = cg_io_outputs_lengths_212; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_213 = cg_io_outputs_lengths_213; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_214 = cg_io_outputs_lengths_214; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_215 = cg_io_outputs_lengths_215; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_216 = cg_io_outputs_lengths_216; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_217 = cg_io_outputs_lengths_217; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_218 = cg_io_outputs_lengths_218; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_219 = cg_io_outputs_lengths_219; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_220 = cg_io_outputs_lengths_220; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_221 = cg_io_outputs_lengths_221; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_222 = cg_io_outputs_lengths_222; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_223 = cg_io_outputs_lengths_223; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_224 = cg_io_outputs_lengths_224; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_225 = cg_io_outputs_lengths_225; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_226 = cg_io_outputs_lengths_226; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_227 = cg_io_outputs_lengths_227; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_228 = cg_io_outputs_lengths_228; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_229 = cg_io_outputs_lengths_229; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_230 = cg_io_outputs_lengths_230; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_231 = cg_io_outputs_lengths_231; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_232 = cg_io_outputs_lengths_232; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_233 = cg_io_outputs_lengths_233; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_234 = cg_io_outputs_lengths_234; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_235 = cg_io_outputs_lengths_235; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_236 = cg_io_outputs_lengths_236; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_237 = cg_io_outputs_lengths_237; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_238 = cg_io_outputs_lengths_238; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_239 = cg_io_outputs_lengths_239; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_240 = cg_io_outputs_lengths_240; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_241 = cg_io_outputs_lengths_241; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_242 = cg_io_outputs_lengths_242; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_243 = cg_io_outputs_lengths_243; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_244 = cg_io_outputs_lengths_244; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_245 = cg_io_outputs_lengths_245; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_246 = cg_io_outputs_lengths_246; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_247 = cg_io_outputs_lengths_247; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_248 = cg_io_outputs_lengths_248; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_249 = cg_io_outputs_lengths_249; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_250 = cg_io_outputs_lengths_250; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_251 = cg_io_outputs_lengths_251; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_252 = cg_io_outputs_lengths_252; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_253 = cg_io_outputs_lengths_253; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_254 = cg_io_outputs_lengths_254; // @[topLevel.scala 102:16]
  assign co_io_inputs_lengths_255 = cg_io_outputs_lengths_255; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_0 = cg_io_outputs_charactersOut_0; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_1 = cg_io_outputs_charactersOut_1; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_2 = cg_io_outputs_charactersOut_2; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_3 = cg_io_outputs_charactersOut_3; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_4 = cg_io_outputs_charactersOut_4; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_5 = cg_io_outputs_charactersOut_5; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_6 = cg_io_outputs_charactersOut_6; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_7 = cg_io_outputs_charactersOut_7; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_8 = cg_io_outputs_charactersOut_8; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_9 = cg_io_outputs_charactersOut_9; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_10 = cg_io_outputs_charactersOut_10; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_11 = cg_io_outputs_charactersOut_11; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_12 = cg_io_outputs_charactersOut_12; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_13 = cg_io_outputs_charactersOut_13; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_14 = cg_io_outputs_charactersOut_14; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_15 = cg_io_outputs_charactersOut_15; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_16 = cg_io_outputs_charactersOut_16; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_17 = cg_io_outputs_charactersOut_17; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_18 = cg_io_outputs_charactersOut_18; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_19 = cg_io_outputs_charactersOut_19; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_20 = cg_io_outputs_charactersOut_20; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_21 = cg_io_outputs_charactersOut_21; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_22 = cg_io_outputs_charactersOut_22; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_23 = cg_io_outputs_charactersOut_23; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_24 = cg_io_outputs_charactersOut_24; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_25 = cg_io_outputs_charactersOut_25; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_26 = cg_io_outputs_charactersOut_26; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_27 = cg_io_outputs_charactersOut_27; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_28 = cg_io_outputs_charactersOut_28; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_29 = cg_io_outputs_charactersOut_29; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_30 = cg_io_outputs_charactersOut_30; // @[topLevel.scala 102:16]
  assign co_io_inputs_charactersOut_31 = cg_io_outputs_charactersOut_31; // @[topLevel.scala 102:16]
  assign co_io_inputs_nodes = cg_io_outputs_nodes; // @[topLevel.scala 102:16]
  assign co_io_inputs_escapeCharacterLength = cg_io_outputs_escapeCharacterLength; // @[topLevel.scala 102:16]
  assign co_io_inputs_escapeCodeword = cg_io_outputs_escapeCodeword; // @[topLevel.scala 102:16]
  assign co_io_outputs_0_ready = io_outputs_0_ready; // @[topLevel.scala 103:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  previousStart = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cfmPreviousFinished = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  tgPreviousFinished = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  tdcPreviousFinished = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  sltgPreviousFinished = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  tnPreviousFinished = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  cgPreviousFinished = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  coPreviousFinished = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    previousStart <= io_start;
    cfmPreviousFinished <= cfm_io_finished;
    tgPreviousFinished <= tg_io_finished;
    tdcPreviousFinished <= tdc_io_finished;
    sltgPreviousFinished <= sltg_io_finished;
    tnPreviousFinished <= tn_io_finished;
    cgPreviousFinished <= cg_io_finished;
    coPreviousFinished <= co_io_finished;
  end
endmodule
module compressorBytesToCacheLine(
  input          clock,
  input          reset,
  output         io_inputData_ready,
  input          io_inputData_valid,
  input  [27:0]  io_inputData_bits,
  input  [4:0]   io_inputDataLength,
  input          io_dumpBuffer,
  output [9:0]   io_currentBufferBits,
  input          io_outputData_ready,
  output         io_outputData_valid,
  output [511:0] io_outputData_bits
);
  reg [9:0] currentBufferBits; // @[compressorBytesToCacheLine.scala 41:34]
  reg [31:0] _RAND_0;
  reg [538:0] buffer; // @[compressorBytesToCacheLine.scala 43:19]
  reg [543:0] _RAND_1;
  wire [538:0] _GEN_1 = io_outputData_ready ? 539'h0 : buffer; // @[compressorBytesToCacheLine.scala 48:31]
  wire  _T = currentBufferBits >= 10'h200; // @[compressorBytesToCacheLine.scala 54:28]
  wire [9:0] _T_2 = currentBufferBits - 10'h200; // @[compressorBytesToCacheLine.scala 60:48]
  wire  _T_3 = currentBufferBits == 10'h200; // @[compressorBytesToCacheLine.scala 61:32]
  wire [1050:0] _T_4 = {buffer, 512'h0}; // @[compressorBytesToCacheLine.scala 64:28]
  wire [1050:0] _GEN_2 = _T_3 ? 1051'h0 : _T_4; // @[compressorBytesToCacheLine.scala 61:54]
  wire [1050:0] _GEN_4 = io_outputData_ready ? _GEN_2 : {{512'd0}, buffer}; // @[compressorBytesToCacheLine.scala 58:33]
  wire [9:0] _GEN_15 = {{5'd0}, io_inputDataLength}; // @[compressorBytesToCacheLine.scala 72:48]
  wire [9:0] _T_6 = currentBufferBits + _GEN_15; // @[compressorBytesToCacheLine.scala 72:48]
  wire [58:0] _T_8 = 59'hfffffff << io_inputDataLength; // @[compressorBytesToCacheLine.scala 73:80]
  wire [58:0] _T_9 = ~_T_8; // @[compressorBytesToCacheLine.scala 73:50]
  wire [58:0] _GEN_16 = {{31'd0}, io_inputData_bits}; // @[compressorBytesToCacheLine.scala 73:48]
  wire [58:0] _T_10 = _GEN_16 & _T_9; // @[compressorBytesToCacheLine.scala 73:48]
  wire [9:0] _T_12 = 10'h21b - _GEN_15; // @[compressorBytesToCacheLine.scala 73:121]
  wire [9:0] _T_14 = _T_12 - currentBufferBits; // @[compressorBytesToCacheLine.scala 73:142]
  wire [1081:0] _GEN_18 = {{1023'd0}, _T_10}; // @[compressorBytesToCacheLine.scala 73:104]
  wire [1081:0] _T_15 = _GEN_18 << _T_14; // @[compressorBytesToCacheLine.scala 73:104]
  wire [1081:0] _GEN_19 = {{543'd0}, buffer}; // @[compressorBytesToCacheLine.scala 73:26]
  wire [1081:0] _T_16 = _GEN_19 | _T_15; // @[compressorBytesToCacheLine.scala 73:26]
  wire [1081:0] _GEN_6 = io_inputData_valid ? _T_16 : {{543'd0}, buffer}; // @[compressorBytesToCacheLine.scala 70:32]
  wire  _GEN_7 = _T ? 1'h0 : 1'h1; // @[compressorBytesToCacheLine.scala 54:49]
  wire [1081:0] _GEN_10 = _T ? {{31'd0}, _GEN_4} : _GEN_6; // @[compressorBytesToCacheLine.scala 54:49]
  wire [1081:0] _GEN_14 = io_dumpBuffer ? {{543'd0}, _GEN_1} : _GEN_10; // @[compressorBytesToCacheLine.scala 45:23]
  assign io_inputData_ready = io_dumpBuffer ? 1'h0 : _GEN_7; // @[compressorBytesToCacheLine.scala 47:24 compressorBytesToCacheLine.scala 56:26 compressorBytesToCacheLine.scala 69:26]
  assign io_currentBufferBits = currentBufferBits; // @[compressorBytesToCacheLine.scala 42:24]
  assign io_outputData_valid = io_dumpBuffer | _T; // @[compressorBytesToCacheLine.scala 46:25 compressorBytesToCacheLine.scala 57:27 compressorBytesToCacheLine.scala 68:27]
  assign io_outputData_bits = buffer[538:27]; // @[compressorBytesToCacheLine.scala 79:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  currentBufferBits = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {17{`RANDOM}};
  buffer = _RAND_1[538:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      currentBufferBits <= 10'h0;
    end else if (io_dumpBuffer) begin
      if (io_outputData_ready) begin
        currentBufferBits <= 10'h0;
      end
    end else if (_T) begin
      if (io_outputData_ready) begin
        currentBufferBits <= _T_2;
      end
    end else if (io_inputData_valid) begin
      currentBufferBits <= _T_6;
    end
    buffer <= _GEN_14[538:0];
  end
endmodule
module huffmanCompressorCacheLineWrapper(
  input          clock,
  input          reset,
  input          io_start,
  output [5:0]   io_readPointer,
  output         io_loadReadPointer,
  input          io_readFifoEmpty,
  output         io_readReady,
  input          io_readValid,
  input  [511:0] io_readData,
  input          io_writeFifoFull,
  output         io_writeRequest,
  output [511:0] io_writeData,
  output [13:0]  io_compressedSize,
  output         io_incompressible,
  output         io_done
);
  reg [7:0] inputDataCache [0:4095]; // @[huffmanCompressorCacheLineWrapper.scala 105:16]
  reg [31:0] _RAND_0;
  wire [7:0] inputDataCache__T_262613_data; // @[huffmanCompressorCacheLineWrapper.scala 105:16]
  wire [11:0] inputDataCache__T_262613_addr; // @[huffmanCompressorCacheLineWrapper.scala 105:16]
  wire [7:0] inputDataCache__T_262608_data; // @[huffmanCompressorCacheLineWrapper.scala 105:16]
  wire [11:0] inputDataCache__T_262608_addr; // @[huffmanCompressorCacheLineWrapper.scala 105:16]
  wire  inputDataCache__T_262608_mask; // @[huffmanCompressorCacheLineWrapper.scala 105:16]
  wire  inputDataCache__T_262608_en; // @[huffmanCompressorCacheLineWrapper.scala 105:16]
  reg  inputDataCache__T_262613_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [11:0] inputDataCache__T_262613_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  compressor_clock; // @[huffmanCompressorCacheLineWrapper.scala 121:26]
  wire  compressor_reset; // @[huffmanCompressorCacheLineWrapper.scala 121:26]
  wire  compressor_io_start; // @[huffmanCompressorCacheLineWrapper.scala 121:26]
  wire [11:0] compressor_io_characterFrequencyInputs_currentByteOut; // @[huffmanCompressorCacheLineWrapper.scala 121:26]
  wire [7:0] compressor_io_characterFrequencyInputs_dataIn_0; // @[huffmanCompressorCacheLineWrapper.scala 121:26]
  wire  compressor_io_characterFrequencyInputs_valid; // @[huffmanCompressorCacheLineWrapper.scala 121:26]
  wire  compressor_io_characterFrequencyInputs_ready; // @[huffmanCompressorCacheLineWrapper.scala 121:26]
  wire [11:0] compressor_io_compressionInputs_0_currentByteOut; // @[huffmanCompressorCacheLineWrapper.scala 121:26]
  wire [7:0] compressor_io_compressionInputs_0_dataIn_0; // @[huffmanCompressorCacheLineWrapper.scala 121:26]
  wire  compressor_io_compressionInputs_0_valid; // @[huffmanCompressorCacheLineWrapper.scala 121:26]
  wire  compressor_io_compressionInputs_0_ready; // @[huffmanCompressorCacheLineWrapper.scala 121:26]
  wire [27:0] compressor_io_outputs_0_dataOut; // @[huffmanCompressorCacheLineWrapper.scala 121:26]
  wire [4:0] compressor_io_outputs_0_dataLength; // @[huffmanCompressorCacheLineWrapper.scala 121:26]
  wire  compressor_io_outputs_0_valid; // @[huffmanCompressorCacheLineWrapper.scala 121:26]
  wire  compressor_io_outputs_0_ready; // @[huffmanCompressorCacheLineWrapper.scala 121:26]
  wire  compressor_io_finished; // @[huffmanCompressorCacheLineWrapper.scala 121:26]
  wire  writeCacheLineConverter_clock; // @[huffmanCompressorCacheLineWrapper.scala 125:39]
  wire  writeCacheLineConverter_reset; // @[huffmanCompressorCacheLineWrapper.scala 125:39]
  wire  writeCacheLineConverter_io_inputData_ready; // @[huffmanCompressorCacheLineWrapper.scala 125:39]
  wire  writeCacheLineConverter_io_inputData_valid; // @[huffmanCompressorCacheLineWrapper.scala 125:39]
  wire [27:0] writeCacheLineConverter_io_inputData_bits; // @[huffmanCompressorCacheLineWrapper.scala 125:39]
  wire [4:0] writeCacheLineConverter_io_inputDataLength; // @[huffmanCompressorCacheLineWrapper.scala 125:39]
  wire  writeCacheLineConverter_io_dumpBuffer; // @[huffmanCompressorCacheLineWrapper.scala 125:39]
  wire [9:0] writeCacheLineConverter_io_currentBufferBits; // @[huffmanCompressorCacheLineWrapper.scala 125:39]
  wire  writeCacheLineConverter_io_outputData_ready; // @[huffmanCompressorCacheLineWrapper.scala 125:39]
  wire  writeCacheLineConverter_io_outputData_valid; // @[huffmanCompressorCacheLineWrapper.scala 125:39]
  wire [511:0] writeCacheLineConverter_io_outputData_bits; // @[huffmanCompressorCacheLineWrapper.scala 125:39]
  wire  readDataAsFlattenedVec_63_0 = io_readData[0]; // @[huffmanCompressorCacheLineWrapper.scala 97:98]
  wire [7:0] readDataAsVec_0 = {io_readData[511],io_readData[510],io_readData[509],io_readData[508],io_readData[507],io_readData[506],io_readData[505],io_readData[504]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_1 = {io_readData[503],io_readData[502],io_readData[501],io_readData[500],io_readData[499],io_readData[498],io_readData[497],io_readData[496]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_2 = {io_readData[495],io_readData[494],io_readData[493],io_readData[492],io_readData[491],io_readData[490],io_readData[489],io_readData[488]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_3 = {io_readData[487],io_readData[486],io_readData[485],io_readData[484],io_readData[483],io_readData[482],io_readData[481],io_readData[480]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_4 = {io_readData[479],io_readData[478],io_readData[477],io_readData[476],io_readData[475],io_readData[474],io_readData[473],io_readData[472]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_5 = {io_readData[471],io_readData[470],io_readData[469],io_readData[468],io_readData[467],io_readData[466],io_readData[465],io_readData[464]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_6 = {io_readData[463],io_readData[462],io_readData[461],io_readData[460],io_readData[459],io_readData[458],io_readData[457],io_readData[456]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_7 = {io_readData[455],io_readData[454],io_readData[453],io_readData[452],io_readData[451],io_readData[450],io_readData[449],io_readData[448]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_8 = {io_readData[447],io_readData[446],io_readData[445],io_readData[444],io_readData[443],io_readData[442],io_readData[441],io_readData[440]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_9 = {io_readData[439],io_readData[438],io_readData[437],io_readData[436],io_readData[435],io_readData[434],io_readData[433],io_readData[432]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_10 = {io_readData[431],io_readData[430],io_readData[429],io_readData[428],io_readData[427],io_readData[426],io_readData[425],io_readData[424]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_11 = {io_readData[423],io_readData[422],io_readData[421],io_readData[420],io_readData[419],io_readData[418],io_readData[417],io_readData[416]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_12 = {io_readData[415],io_readData[414],io_readData[413],io_readData[412],io_readData[411],io_readData[410],io_readData[409],io_readData[408]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_13 = {io_readData[407],io_readData[406],io_readData[405],io_readData[404],io_readData[403],io_readData[402],io_readData[401],io_readData[400]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_14 = {io_readData[399],io_readData[398],io_readData[397],io_readData[396],io_readData[395],io_readData[394],io_readData[393],io_readData[392]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_15 = {io_readData[391],io_readData[390],io_readData[389],io_readData[388],io_readData[387],io_readData[386],io_readData[385],io_readData[384]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_16 = {io_readData[383],io_readData[382],io_readData[381],io_readData[380],io_readData[379],io_readData[378],io_readData[377],io_readData[376]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_17 = {io_readData[375],io_readData[374],io_readData[373],io_readData[372],io_readData[371],io_readData[370],io_readData[369],io_readData[368]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_18 = {io_readData[367],io_readData[366],io_readData[365],io_readData[364],io_readData[363],io_readData[362],io_readData[361],io_readData[360]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_19 = {io_readData[359],io_readData[358],io_readData[357],io_readData[356],io_readData[355],io_readData[354],io_readData[353],io_readData[352]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_20 = {io_readData[351],io_readData[350],io_readData[349],io_readData[348],io_readData[347],io_readData[346],io_readData[345],io_readData[344]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_21 = {io_readData[343],io_readData[342],io_readData[341],io_readData[340],io_readData[339],io_readData[338],io_readData[337],io_readData[336]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_22 = {io_readData[335],io_readData[334],io_readData[333],io_readData[332],io_readData[331],io_readData[330],io_readData[329],io_readData[328]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_23 = {io_readData[327],io_readData[326],io_readData[325],io_readData[324],io_readData[323],io_readData[322],io_readData[321],io_readData[320]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_24 = {io_readData[319],io_readData[318],io_readData[317],io_readData[316],io_readData[315],io_readData[314],io_readData[313],io_readData[312]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_25 = {io_readData[311],io_readData[310],io_readData[309],io_readData[308],io_readData[307],io_readData[306],io_readData[305],io_readData[304]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_26 = {io_readData[303],io_readData[302],io_readData[301],io_readData[300],io_readData[299],io_readData[298],io_readData[297],io_readData[296]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_27 = {io_readData[295],io_readData[294],io_readData[293],io_readData[292],io_readData[291],io_readData[290],io_readData[289],io_readData[288]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_28 = {io_readData[287],io_readData[286],io_readData[285],io_readData[284],io_readData[283],io_readData[282],io_readData[281],io_readData[280]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_29 = {io_readData[279],io_readData[278],io_readData[277],io_readData[276],io_readData[275],io_readData[274],io_readData[273],io_readData[272]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_30 = {io_readData[271],io_readData[270],io_readData[269],io_readData[268],io_readData[267],io_readData[266],io_readData[265],io_readData[264]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_31 = {io_readData[263],io_readData[262],io_readData[261],io_readData[260],io_readData[259],io_readData[258],io_readData[257],io_readData[256]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_32 = {io_readData[255],io_readData[254],io_readData[253],io_readData[252],io_readData[251],io_readData[250],io_readData[249],io_readData[248]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_33 = {io_readData[247],io_readData[246],io_readData[245],io_readData[244],io_readData[243],io_readData[242],io_readData[241],io_readData[240]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_34 = {io_readData[239],io_readData[238],io_readData[237],io_readData[236],io_readData[235],io_readData[234],io_readData[233],io_readData[232]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_35 = {io_readData[231],io_readData[230],io_readData[229],io_readData[228],io_readData[227],io_readData[226],io_readData[225],io_readData[224]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_36 = {io_readData[223],io_readData[222],io_readData[221],io_readData[220],io_readData[219],io_readData[218],io_readData[217],io_readData[216]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_37 = {io_readData[215],io_readData[214],io_readData[213],io_readData[212],io_readData[211],io_readData[210],io_readData[209],io_readData[208]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_38 = {io_readData[207],io_readData[206],io_readData[205],io_readData[204],io_readData[203],io_readData[202],io_readData[201],io_readData[200]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_39 = {io_readData[199],io_readData[198],io_readData[197],io_readData[196],io_readData[195],io_readData[194],io_readData[193],io_readData[192]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_40 = {io_readData[191],io_readData[190],io_readData[189],io_readData[188],io_readData[187],io_readData[186],io_readData[185],io_readData[184]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_41 = {io_readData[183],io_readData[182],io_readData[181],io_readData[180],io_readData[179],io_readData[178],io_readData[177],io_readData[176]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_42 = {io_readData[175],io_readData[174],io_readData[173],io_readData[172],io_readData[171],io_readData[170],io_readData[169],io_readData[168]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_43 = {io_readData[167],io_readData[166],io_readData[165],io_readData[164],io_readData[163],io_readData[162],io_readData[161],io_readData[160]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_44 = {io_readData[159],io_readData[158],io_readData[157],io_readData[156],io_readData[155],io_readData[154],io_readData[153],io_readData[152]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_45 = {io_readData[151],io_readData[150],io_readData[149],io_readData[148],io_readData[147],io_readData[146],io_readData[145],io_readData[144]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_46 = {io_readData[143],io_readData[142],io_readData[141],io_readData[140],io_readData[139],io_readData[138],io_readData[137],io_readData[136]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_47 = {io_readData[135],io_readData[134],io_readData[133],io_readData[132],io_readData[131],io_readData[130],io_readData[129],io_readData[128]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_48 = {io_readData[127],io_readData[126],io_readData[125],io_readData[124],io_readData[123],io_readData[122],io_readData[121],io_readData[120]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_49 = {io_readData[119],io_readData[118],io_readData[117],io_readData[116],io_readData[115],io_readData[114],io_readData[113],io_readData[112]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_50 = {io_readData[111],io_readData[110],io_readData[109],io_readData[108],io_readData[107],io_readData[106],io_readData[105],io_readData[104]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_51 = {io_readData[103],io_readData[102],io_readData[101],io_readData[100],io_readData[99],io_readData[98],io_readData[97],io_readData[96]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_52 = {io_readData[95],io_readData[94],io_readData[93],io_readData[92],io_readData[91],io_readData[90],io_readData[89],io_readData[88]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_53 = {io_readData[87],io_readData[86],io_readData[85],io_readData[84],io_readData[83],io_readData[82],io_readData[81],io_readData[80]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_54 = {io_readData[79],io_readData[78],io_readData[77],io_readData[76],io_readData[75],io_readData[74],io_readData[73],io_readData[72]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_55 = {io_readData[71],io_readData[70],io_readData[69],io_readData[68],io_readData[67],io_readData[66],io_readData[65],io_readData[64]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_56 = {io_readData[63],io_readData[62],io_readData[61],io_readData[60],io_readData[59],io_readData[58],io_readData[57],io_readData[56]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_57 = {io_readData[55],io_readData[54],io_readData[53],io_readData[52],io_readData[51],io_readData[50],io_readData[49],io_readData[48]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_58 = {io_readData[47],io_readData[46],io_readData[45],io_readData[44],io_readData[43],io_readData[42],io_readData[41],io_readData[40]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_59 = {io_readData[39],io_readData[38],io_readData[37],io_readData[36],io_readData[35],io_readData[34],io_readData[33],io_readData[32]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_60 = {io_readData[31],io_readData[30],io_readData[29],io_readData[28],io_readData[27],io_readData[26],io_readData[25],io_readData[24]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_61 = {io_readData[23],io_readData[22],io_readData[21],io_readData[20],io_readData[19],io_readData[18],io_readData[17],io_readData[16]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_62 = {io_readData[15],io_readData[14],io_readData[13],io_readData[12],io_readData[11],io_readData[10],io_readData[9],io_readData[8]}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  wire [7:0] readDataAsVec_63 = {io_readData[7],io_readData[6],io_readData[5],io_readData[4],io_readData[3],io_readData[2],io_readData[1],readDataAsFlattenedVec_63_0}; // @[huffmanCompressorCacheLineWrapper.scala 99:75]
  reg [7:0] inputDataCacheByte; // @[huffmanCompressorCacheLineWrapper.scala 107:31]
  reg [31:0] _RAND_3;
  reg [2:0] state; // @[huffmanCompressorCacheLineWrapper.scala 114:22]
  reg [31:0] _RAND_4;
  reg [6:0] iterations; // @[huffmanCompressorCacheLineWrapper.scala 116:27]
  reg [31:0] _RAND_5;
  reg [13:0] compressedSize; // @[huffmanCompressorCacheLineWrapper.scala 119:31]
  reg [31:0] _RAND_6;
  wire  _T_262592 = state == 3'h5; // @[huffmanCompressorCacheLineWrapper.scala 138:20]
  wire  _T_262593 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_262594 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire [11:0] _T_262595 = compressor_io_characterFrequencyInputs_currentByteOut / 12'h40; // @[huffmanCompressorCacheLineWrapper.scala 167:79]
  wire  _T_262596 = ~compressor_io_compressionInputs_0_ready; // @[huffmanCompressorCacheLineWrapper.scala 168:12]
  wire  _GEN_3 = compressor_io_characterFrequencyInputs_ready & io_readFifoEmpty; // @[huffmanCompressorCacheLineWrapper.scala 169:60]
  wire  _GEN_5 = _T_262596 & _GEN_3; // @[huffmanCompressorCacheLineWrapper.scala 168:55]
  wire  _T_262597 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_262598 = iterations >= 7'h40; // @[huffmanCompressorCacheLineWrapper.scala 184:25]
  wire [6:0] _T_262600 = iterations + 7'h1; // @[huffmanCompressorCacheLineWrapper.scala 193:38]
  wire [7:0] _T_262601 = iterations * 7'h1; // @[huffmanCompressorCacheLineWrapper.scala 195:56]
  wire [8:0] _T_262602 = {{1'd0}, _T_262601}; // @[huffmanCompressorCacheLineWrapper.scala 195:43]
  wire [12:0] _T_262604 = {{1'd0}, compressor_io_characterFrequencyInputs_currentByteOut}; // @[huffmanCompressorCacheLineWrapper.scala 196:95]
  wire [7:0] _GEN_8 = 6'h1 == _T_262602[5:0] ? readDataAsVec_1 : readDataAsVec_0; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_9 = 6'h2 == _T_262602[5:0] ? readDataAsVec_2 : _GEN_8; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_10 = 6'h3 == _T_262602[5:0] ? readDataAsVec_3 : _GEN_9; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_11 = 6'h4 == _T_262602[5:0] ? readDataAsVec_4 : _GEN_10; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_12 = 6'h5 == _T_262602[5:0] ? readDataAsVec_5 : _GEN_11; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_13 = 6'h6 == _T_262602[5:0] ? readDataAsVec_6 : _GEN_12; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_14 = 6'h7 == _T_262602[5:0] ? readDataAsVec_7 : _GEN_13; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_15 = 6'h8 == _T_262602[5:0] ? readDataAsVec_8 : _GEN_14; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_16 = 6'h9 == _T_262602[5:0] ? readDataAsVec_9 : _GEN_15; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_17 = 6'ha == _T_262602[5:0] ? readDataAsVec_10 : _GEN_16; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_18 = 6'hb == _T_262602[5:0] ? readDataAsVec_11 : _GEN_17; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_19 = 6'hc == _T_262602[5:0] ? readDataAsVec_12 : _GEN_18; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_20 = 6'hd == _T_262602[5:0] ? readDataAsVec_13 : _GEN_19; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_21 = 6'he == _T_262602[5:0] ? readDataAsVec_14 : _GEN_20; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_22 = 6'hf == _T_262602[5:0] ? readDataAsVec_15 : _GEN_21; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_23 = 6'h10 == _T_262602[5:0] ? readDataAsVec_16 : _GEN_22; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_24 = 6'h11 == _T_262602[5:0] ? readDataAsVec_17 : _GEN_23; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_25 = 6'h12 == _T_262602[5:0] ? readDataAsVec_18 : _GEN_24; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_26 = 6'h13 == _T_262602[5:0] ? readDataAsVec_19 : _GEN_25; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_27 = 6'h14 == _T_262602[5:0] ? readDataAsVec_20 : _GEN_26; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_28 = 6'h15 == _T_262602[5:0] ? readDataAsVec_21 : _GEN_27; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_29 = 6'h16 == _T_262602[5:0] ? readDataAsVec_22 : _GEN_28; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_30 = 6'h17 == _T_262602[5:0] ? readDataAsVec_23 : _GEN_29; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_31 = 6'h18 == _T_262602[5:0] ? readDataAsVec_24 : _GEN_30; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_32 = 6'h19 == _T_262602[5:0] ? readDataAsVec_25 : _GEN_31; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_33 = 6'h1a == _T_262602[5:0] ? readDataAsVec_26 : _GEN_32; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_34 = 6'h1b == _T_262602[5:0] ? readDataAsVec_27 : _GEN_33; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_35 = 6'h1c == _T_262602[5:0] ? readDataAsVec_28 : _GEN_34; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_36 = 6'h1d == _T_262602[5:0] ? readDataAsVec_29 : _GEN_35; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_37 = 6'h1e == _T_262602[5:0] ? readDataAsVec_30 : _GEN_36; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_38 = 6'h1f == _T_262602[5:0] ? readDataAsVec_31 : _GEN_37; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_39 = 6'h20 == _T_262602[5:0] ? readDataAsVec_32 : _GEN_38; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_40 = 6'h21 == _T_262602[5:0] ? readDataAsVec_33 : _GEN_39; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_41 = 6'h22 == _T_262602[5:0] ? readDataAsVec_34 : _GEN_40; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_42 = 6'h23 == _T_262602[5:0] ? readDataAsVec_35 : _GEN_41; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_43 = 6'h24 == _T_262602[5:0] ? readDataAsVec_36 : _GEN_42; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_44 = 6'h25 == _T_262602[5:0] ? readDataAsVec_37 : _GEN_43; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_45 = 6'h26 == _T_262602[5:0] ? readDataAsVec_38 : _GEN_44; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_46 = 6'h27 == _T_262602[5:0] ? readDataAsVec_39 : _GEN_45; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_47 = 6'h28 == _T_262602[5:0] ? readDataAsVec_40 : _GEN_46; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_48 = 6'h29 == _T_262602[5:0] ? readDataAsVec_41 : _GEN_47; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_49 = 6'h2a == _T_262602[5:0] ? readDataAsVec_42 : _GEN_48; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_50 = 6'h2b == _T_262602[5:0] ? readDataAsVec_43 : _GEN_49; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_51 = 6'h2c == _T_262602[5:0] ? readDataAsVec_44 : _GEN_50; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_52 = 6'h2d == _T_262602[5:0] ? readDataAsVec_45 : _GEN_51; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_53 = 6'h2e == _T_262602[5:0] ? readDataAsVec_46 : _GEN_52; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_54 = 6'h2f == _T_262602[5:0] ? readDataAsVec_47 : _GEN_53; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_55 = 6'h30 == _T_262602[5:0] ? readDataAsVec_48 : _GEN_54; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_56 = 6'h31 == _T_262602[5:0] ? readDataAsVec_49 : _GEN_55; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_57 = 6'h32 == _T_262602[5:0] ? readDataAsVec_50 : _GEN_56; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_58 = 6'h33 == _T_262602[5:0] ? readDataAsVec_51 : _GEN_57; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_59 = 6'h34 == _T_262602[5:0] ? readDataAsVec_52 : _GEN_58; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_60 = 6'h35 == _T_262602[5:0] ? readDataAsVec_53 : _GEN_59; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_61 = 6'h36 == _T_262602[5:0] ? readDataAsVec_54 : _GEN_60; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_62 = 6'h37 == _T_262602[5:0] ? readDataAsVec_55 : _GEN_61; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_63 = 6'h38 == _T_262602[5:0] ? readDataAsVec_56 : _GEN_62; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_64 = 6'h39 == _T_262602[5:0] ? readDataAsVec_57 : _GEN_63; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_65 = 6'h3a == _T_262602[5:0] ? readDataAsVec_58 : _GEN_64; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_66 = 6'h3b == _T_262602[5:0] ? readDataAsVec_59 : _GEN_65; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_67 = 6'h3c == _T_262602[5:0] ? readDataAsVec_60 : _GEN_66; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_68 = 6'h3d == _T_262602[5:0] ? readDataAsVec_61 : _GEN_67; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_69 = 6'h3e == _T_262602[5:0] ? readDataAsVec_62 : _GEN_68; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_70 = 6'h3f == _T_262602[5:0] ? readDataAsVec_63 : _GEN_69; // @[huffmanCompressorCacheLineWrapper.scala 197:68]
  wire [7:0] _GEN_136 = compressor_io_characterFrequencyInputs_ready ? _GEN_70 : 8'h0; // @[huffmanCompressorCacheLineWrapper.scala 190:62]
  wire  _GEN_139 = compressor_io_characterFrequencyInputs_ready; // @[huffmanCompressorCacheLineWrapper.scala 190:62]
  wire  _GEN_144 = _T_262598 ? 1'h0 : 1'h1; // @[huffmanCompressorCacheLineWrapper.scala 184:56]
  wire [7:0] _GEN_146 = _T_262598 ? 8'h0 : _GEN_136; // @[huffmanCompressorCacheLineWrapper.scala 184:56]
  wire  _GEN_149 = _T_262598 ? 1'h0 : _GEN_139; // @[huffmanCompressorCacheLineWrapper.scala 184:56]
  wire  _GEN_153 = io_readValid & _T_262598; // @[huffmanCompressorCacheLineWrapper.scala 182:26]
  wire  _GEN_154 = io_readValid & _GEN_144; // @[huffmanCompressorCacheLineWrapper.scala 182:26]
  wire [7:0] _GEN_156 = io_readValid ? _GEN_146 : 8'h0; // @[huffmanCompressorCacheLineWrapper.scala 182:26]
  wire  _GEN_159 = io_readValid & _GEN_149; // @[huffmanCompressorCacheLineWrapper.scala 182:26]
  wire  _T_262609 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_262610 = writeCacheLineConverter_io_currentBufferBits > 10'h0; // @[huffmanCompressorCacheLineWrapper.scala 208:59]
  wire  _T_262611 = ~io_writeFifoFull; // @[huffmanCompressorCacheLineWrapper.scala 212:18]
  wire  _GEN_163 = writeCacheLineConverter_io_outputData_valid & _T_262611; // @[huffmanCompressorCacheLineWrapper.scala 211:61]
  wire  _GEN_165 = _T_262610 & _GEN_163; // @[huffmanCompressorCacheLineWrapper.scala 208:66]
  wire  _GEN_170 = compressor_io_compressionInputs_0_ready; // @[huffmanCompressorCacheLineWrapper.scala 229:58]
  wire  _GEN_176 = writeCacheLineConverter_io_outputData_valid ? 1'h0 : _GEN_170; // @[huffmanCompressorCacheLineWrapper.scala 222:59]
  wire  _GEN_179 = compressor_io_finished & _T_262610; // @[huffmanCompressorCacheLineWrapper.scala 206:36]
  wire  _GEN_180 = compressor_io_finished ? _GEN_165 : _GEN_163; // @[huffmanCompressorCacheLineWrapper.scala 206:36]
  wire  _GEN_184 = compressor_io_finished ? 1'h0 : _GEN_176; // @[huffmanCompressorCacheLineWrapper.scala 206:36]
  wire  _T_262614 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_262615 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_262616 = ~io_start; // @[huffmanCompressorCacheLineWrapper.scala 246:12]
  wire  _GEN_188 = _T_262615 | _T_262592; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_191 = _T_262614 ? inputDataCacheByte : 8'h0; // @[Conditional.scala 39:67]
  wire  _GEN_193 = _T_262614 ? _T_262592 : _GEN_188; // @[Conditional.scala 39:67]
  wire  _GEN_194 = _T_262609 & _GEN_179; // @[Conditional.scala 39:67]
  wire  _GEN_195 = _T_262609 & _GEN_180; // @[Conditional.scala 39:67]
  wire  _GEN_199 = _T_262609 & _GEN_184; // @[Conditional.scala 39:67]
  wire  _GEN_201 = _T_262609 ? 1'h0 : _T_262614; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_202 = _T_262609 ? 8'h0 : _GEN_191; // @[Conditional.scala 39:67]
  wire  _GEN_203 = _T_262609 ? _T_262592 : _GEN_193; // @[Conditional.scala 39:67]
  wire  _GEN_205 = _T_262597 & _GEN_153; // @[Conditional.scala 39:67]
  wire  _GEN_206 = _T_262597 & _GEN_154; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_208 = _T_262597 ? _GEN_156 : 8'h0; // @[Conditional.scala 39:67]
  wire  _GEN_211 = _T_262597 & _GEN_159; // @[Conditional.scala 39:67]
  wire  _GEN_214 = _T_262597 ? 1'h0 : _GEN_194; // @[Conditional.scala 39:67]
  wire  _GEN_215 = _T_262597 ? 1'h0 : _GEN_195; // @[Conditional.scala 39:67]
  wire  _GEN_218 = _T_262597 ? 1'h0 : _GEN_199; // @[Conditional.scala 39:67]
  wire  _GEN_220 = _T_262597 ? 1'h0 : _GEN_201; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_221 = _T_262597 ? 8'h0 : _GEN_202; // @[Conditional.scala 39:67]
  wire  _GEN_222 = _T_262597 ? _T_262592 : _GEN_203; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_224 = _T_262594 ? _T_262595 : 12'h0; // @[Conditional.scala 39:67]
  wire  _GEN_225 = _T_262594 & _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_227 = _T_262594 ? 1'h0 : _GEN_205; // @[Conditional.scala 39:67]
  wire  _GEN_228 = _T_262594 ? 1'h0 : _GEN_206; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_229 = _T_262594 ? 8'h0 : _GEN_208; // @[Conditional.scala 39:67]
  wire  _GEN_232 = _T_262594 ? 1'h0 : _GEN_211; // @[Conditional.scala 39:67]
  wire  _GEN_235 = _T_262594 ? 1'h0 : _GEN_214; // @[Conditional.scala 39:67]
  wire  _GEN_236 = _T_262594 ? 1'h0 : _GEN_215; // @[Conditional.scala 39:67]
  wire  _GEN_239 = _T_262594 ? 1'h0 : _GEN_218; // @[Conditional.scala 39:67]
  wire  _GEN_241 = _T_262594 ? 1'h0 : _GEN_220; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_242 = _T_262594 ? 8'h0 : _GEN_221; // @[Conditional.scala 39:67]
  wire  _GEN_243 = _T_262594 ? _T_262592 : _GEN_222; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_247 = _T_262593 ? 12'h0 : _GEN_224; // @[Conditional.scala 40:58]
  wire [13:0] _T_262618 = compressedSize + 14'h40; // @[huffmanCompressorCacheLineWrapper.scala 253:38]
  topLevel compressor ( // @[huffmanCompressorCacheLineWrapper.scala 121:26]
    .clock(compressor_clock),
    .reset(compressor_reset),
    .io_start(compressor_io_start),
    .io_characterFrequencyInputs_currentByteOut(compressor_io_characterFrequencyInputs_currentByteOut),
    .io_characterFrequencyInputs_dataIn_0(compressor_io_characterFrequencyInputs_dataIn_0),
    .io_characterFrequencyInputs_valid(compressor_io_characterFrequencyInputs_valid),
    .io_characterFrequencyInputs_ready(compressor_io_characterFrequencyInputs_ready),
    .io_compressionInputs_0_currentByteOut(compressor_io_compressionInputs_0_currentByteOut),
    .io_compressionInputs_0_dataIn_0(compressor_io_compressionInputs_0_dataIn_0),
    .io_compressionInputs_0_valid(compressor_io_compressionInputs_0_valid),
    .io_compressionInputs_0_ready(compressor_io_compressionInputs_0_ready),
    .io_outputs_0_dataOut(compressor_io_outputs_0_dataOut),
    .io_outputs_0_dataLength(compressor_io_outputs_0_dataLength),
    .io_outputs_0_valid(compressor_io_outputs_0_valid),
    .io_outputs_0_ready(compressor_io_outputs_0_ready),
    .io_finished(compressor_io_finished)
  );
  compressorBytesToCacheLine writeCacheLineConverter ( // @[huffmanCompressorCacheLineWrapper.scala 125:39]
    .clock(writeCacheLineConverter_clock),
    .reset(writeCacheLineConverter_reset),
    .io_inputData_ready(writeCacheLineConverter_io_inputData_ready),
    .io_inputData_valid(writeCacheLineConverter_io_inputData_valid),
    .io_inputData_bits(writeCacheLineConverter_io_inputData_bits),
    .io_inputDataLength(writeCacheLineConverter_io_inputDataLength),
    .io_dumpBuffer(writeCacheLineConverter_io_dumpBuffer),
    .io_currentBufferBits(writeCacheLineConverter_io_currentBufferBits),
    .io_outputData_ready(writeCacheLineConverter_io_outputData_ready),
    .io_outputData_valid(writeCacheLineConverter_io_outputData_valid),
    .io_outputData_bits(writeCacheLineConverter_io_outputData_bits)
  );
  assign inputDataCache__T_262613_addr = inputDataCache__T_262613_addr_pipe_0;
  assign inputDataCache__T_262613_data = inputDataCache[inputDataCache__T_262613_addr]; // @[huffmanCompressorCacheLineWrapper.scala 105:16]
  assign inputDataCache__T_262608_data = 6'h3f == _T_262602[5:0] ? readDataAsVec_63 : _GEN_69;
  assign inputDataCache__T_262608_addr = _T_262604[11:0];
  assign inputDataCache__T_262608_mask = 1'h1;
  assign inputDataCache__T_262608_en = _T_262593 ? 1'h0 : _GEN_232;
  assign io_readPointer = _GEN_247[5:0]; // @[huffmanCompressorCacheLineWrapper.scala 146:18 huffmanCompressorCacheLineWrapper.scala 167:22]
  assign io_loadReadPointer = _T_262593 ? 1'h0 : _GEN_225; // @[huffmanCompressorCacheLineWrapper.scala 147:22 huffmanCompressorCacheLineWrapper.scala 172:32]
  assign io_readReady = _T_262593 ? 1'h0 : _GEN_227; // @[huffmanCompressorCacheLineWrapper.scala 145:16 huffmanCompressorCacheLineWrapper.scala 187:24]
  assign io_writeRequest = _T_262593 ? 1'h0 : _GEN_236; // @[huffmanCompressorCacheLineWrapper.scala 150:19 huffmanCompressorCacheLineWrapper.scala 214:31 huffmanCompressorCacheLineWrapper.scala 226:29]
  assign io_writeData = writeCacheLineConverter_io_outputData_bits; // @[huffmanCompressorCacheLineWrapper.scala 132:46]
  assign io_compressedSize = compressedSize; // @[huffmanCompressorCacheLineWrapper.scala 139:21]
  assign io_incompressible = 1'h0; // @[huffmanCompressorCacheLineWrapper.scala 142:21]
  assign io_done = _T_262593 ? _T_262592 : _GEN_243; // @[huffmanCompressorCacheLineWrapper.scala 138:11 huffmanCompressorCacheLineWrapper.scala 245:15]
  assign compressor_clock = clock;
  assign compressor_reset = reset;
  assign compressor_io_start = io_start; // @[huffmanCompressorCacheLineWrapper.scala 122:23]
  assign compressor_io_characterFrequencyInputs_dataIn_0 = _T_262593 ? 8'h0 : _GEN_229; // @[huffmanCompressorCacheLineWrapper.scala 155:58 huffmanCompressorCacheLineWrapper.scala 197:68]
  assign compressor_io_characterFrequencyInputs_valid = _T_262593 ? 1'h0 : _GEN_228; // @[huffmanCompressorCacheLineWrapper.scala 151:48 huffmanCompressorCacheLineWrapper.scala 189:56]
  assign compressor_io_compressionInputs_0_dataIn_0 = _T_262593 ? 8'h0 : _GEN_242; // @[huffmanCompressorCacheLineWrapper.scala 152:48 huffmanCompressorCacheLineWrapper.scala 239:52]
  assign compressor_io_compressionInputs_0_valid = _T_262593 ? 1'h0 : _GEN_241; // @[huffmanCompressorCacheLineWrapper.scala 153:44 huffmanCompressorCacheLineWrapper.scala 238:48]
  assign compressor_io_outputs_0_ready = writeCacheLineConverter_io_inputData_ready; // @[huffmanCompressorCacheLineWrapper.scala 134:46]
  assign writeCacheLineConverter_clock = clock;
  assign writeCacheLineConverter_reset = reset;
  assign writeCacheLineConverter_io_inputData_valid = compressor_io_outputs_0_valid; // @[huffmanCompressorCacheLineWrapper.scala 135:46]
  assign writeCacheLineConverter_io_inputData_bits = compressor_io_outputs_0_dataOut; // @[huffmanCompressorCacheLineWrapper.scala 133:45]
  assign writeCacheLineConverter_io_inputDataLength = compressor_io_outputs_0_dataLength; // @[huffmanCompressorCacheLineWrapper.scala 136:46]
  assign writeCacheLineConverter_io_dumpBuffer = _T_262593 ? 1'h0 : _GEN_235; // @[huffmanCompressorCacheLineWrapper.scala 149:41 huffmanCompressorCacheLineWrapper.scala 210:49]
  assign writeCacheLineConverter_io_outputData_ready = _T_262593 ? 1'h0 : _GEN_236; // @[huffmanCompressorCacheLineWrapper.scala 148:47 huffmanCompressorCacheLineWrapper.scala 213:59 huffmanCompressorCacheLineWrapper.scala 225:57]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4096; initvar = initvar+1)
    inputDataCache[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  inputDataCache__T_262613_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  inputDataCache__T_262613_addr_pipe_0 = _RAND_2[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  inputDataCacheByte = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  iterations = _RAND_5[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  compressedSize = _RAND_6[13:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(inputDataCache__T_262608_en & inputDataCache__T_262608_mask) begin
      inputDataCache[inputDataCache__T_262608_addr] <= inputDataCache__T_262608_data; // @[huffmanCompressorCacheLineWrapper.scala 105:16]
    end
    if (_T_262593) begin
      inputDataCache__T_262613_en_pipe_0 <= 1'h0;
    end else if (_T_262594) begin
      inputDataCache__T_262613_en_pipe_0 <= 1'h0;
    end else if (_T_262597) begin
      inputDataCache__T_262613_en_pipe_0 <= 1'h0;
    end else begin
      inputDataCache__T_262613_en_pipe_0 <= _GEN_199;
    end
    if (_T_262593 ? 1'h0 : _GEN_239) begin
      inputDataCache__T_262613_addr_pipe_0 <= compressor_io_compressionInputs_0_currentByteOut;
    end
    if (!(_T_262593)) begin
      if (!(_T_262594)) begin
        if (!(_T_262597)) begin
          if (_T_262609) begin
            if (!(compressor_io_finished)) begin
              if (!(writeCacheLineConverter_io_outputData_valid)) begin
                if (compressor_io_compressionInputs_0_ready) begin
                  inputDataCacheByte <= inputDataCache__T_262613_data;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 3'h0;
    end else if (_T_262593) begin
      if (io_start) begin
        state <= 3'h1;
      end
    end else if (_T_262594) begin
      if (_T_262596) begin
        if (compressor_io_characterFrequencyInputs_ready) begin
          if (io_readFifoEmpty) begin
            state <= 3'h2;
          end
        end
      end else begin
        state <= 3'h3;
      end
    end else if (_T_262597) begin
      if (io_readValid) begin
        if (_T_262598) begin
          state <= 3'h1;
        end
      end
    end else if (_T_262609) begin
      if (compressor_io_finished) begin
        if (!(_T_262610)) begin
          state <= 3'h5;
        end
      end else if (!(writeCacheLineConverter_io_outputData_valid)) begin
        if (compressor_io_compressionInputs_0_ready) begin
          state <= 3'h4;
        end
      end
    end else if (_T_262614) begin
      if (compressor_io_compressionInputs_0_ready) begin
        state <= 3'h3;
      end
    end else if (_T_262615) begin
      if (_T_262616) begin
        state <= 3'h0;
      end
    end
    if (reset) begin
      iterations <= 7'h0;
    end else if (!(_T_262593)) begin
      if (_T_262594) begin
        iterations <= 7'h0;
      end else if (_T_262597) begin
        if (io_readValid) begin
          if (!(_T_262598)) begin
            if (compressor_io_characterFrequencyInputs_ready) begin
              iterations <= _T_262600;
            end
          end
        end
      end
    end
    if (reset) begin
      compressedSize <= 14'h0;
    end else if (io_writeRequest) begin
      compressedSize <= _T_262618;
    end else if (_T_262593) begin
      compressedSize <= 14'h0;
    end
  end
endmodule
