/////////////////////////////////////////////////////////////////////////////////
//
// Heap Lab Research
// Block : Hawk Control Unit 
// 
// Author : Raghavendra Srinivas
// Contact : raghavs@vt.edu	
/////////////////////////////////////////////////////////////////////////////////
// Description: Unit to control and manage entire hawk operations.
// 		Architecture plan is to pipeline multiple requests of CPU, and
// 		this unit take care off look up att table (with local att cache as
// 		planned in previous architecture) , find victim page to
// 		compress, or uncompress compressed page. Deliver this
// 		compress/uncompress burst mode to read and write page
// 		managers, while control unit can paralley lookup for pending
// 		requests.
// 		But for bringup, this majority of operations is handled by page
// 		managers itself.
// 		So, control unit here is really light now
/////////////////////////////////////////////////////////////////////////////////
//local defines
`define FSM_WID 4
module hawk_ctrl_unit #()
(

    input clk_i,
    input rst_ni,

    //pg_writer handshake
    input init_att_done,
    input init_list_done,
    input tbl_update_done,

    //pg_rdmanager
    input pgrd_mngr_ready,
    input allow_cpu_access,
    input tbl_update,
    
    //cpu master handshake
    output hacd_pkg::cpu_rd_reqpkt_t cpu_rd_reqpkt, 
    output hacd_pkg::cpu_wr_reqpkt_t cpu_wr_reqpkt, 
     
    //to control with hawk_pg_writer
    output logic init_att,
    output logic init_list,
    
    //to control cpu interface
    output logic allow_cpu_rd_access,
    output logic allow_cpu_wr_access
);



//local variables
att_lkup_reqpkt_t lkup_reqpkt,n_lkup_reqpkt;
logic n_allow_cpu_wr_access, n_allow_cpu_rd_access;
logic n_init_att,n_init_list;
logic [`FSM_WID-1:0] n_state;
logic [`FSM_WID-1:0] p_state;
//states
localparam IDLE			='d0,
	   CHK_RD_ACTIVE 	='d1,
	   CHK_WR_ACTIVE 	='d2,
	   RD_LOOKUP_ALLOCATE	='d3,
	   WR_LOOKUP_ALLOCATE	='d4,
	   RD_TBL_UPDATE	='d5,
	   WR_TBL_UPDATE	='d6;

//state & output register
always_ff@(posedge clk_i or negedge rst_ni) 
begin
	if(!rst_ni) begin
		p_state<=IDLE;

		//output regs
		init_att<=1'b1; //init_att is enabled upon reset
		init_list<=1'b1; //init_att is enabled upon reset
	end
	else begin
		p_state<=n_state;

		//output regs
		init_att<=n_init_att;
		init_list<=n_init_list;
	end
end

//fsm combo
always_comb
begin
	n_state=p_state;
	n_init_att=init_att;
	n_init_list=init_list;
	n_allow_cpu_wr_access=0;
	n_allow_cpu_rd_access=0;
	n_lkup_reqpkt='d0;
	case(p_state)
		IDLE: begin
			if(init_att_done) begin //wait in same state till table initialiation is done
				n_init_att=1'b0;
			end
			else if (init_list_done) begin
				n_init_list=1'b0;
				n_state=CHK_RD_ACTIVE;
			end
		end
		CHK_RD_ACTIVE:begin
			if(pgrd_mngr_ready && !allow_cpu_rd_access) begin
				if      (cpu_rd_reqpkt.valid) begin 
					n_lkup_reqpkt.lookup=1'b1;
					n_lkup_reqpkt.hppa=cpu_rd_reqpkt.hppa;	 
				  	n_state=RD_LOOKUP_ALLOCATE;
				end
				else if (cpu_wr_reqpkt.valid) begin
					n_lkup_reqpkt.lookup=1'b1;
					n_lkup_reqpkt.hppa=cpu_wr_reqpkt.hppa;	 
				  	n_state=WR_LOOKUP_ALLOCATE;
		  		end
			end 
			//chk if we need fairness among wries and read later
			//however even if we priotise reads over
			//writes, coherecny should not be breoken, even if read
			//comes on same line as write, which is not yet written. It
			//should be handled at system level /one cache before memory
			//controller
		end
		CHK_WR_ACTIVE: begin
			if(pgrd_mngr_ready && !allow_cpu_wr_access) begin
			       if 	(cpu_wr_reqpkt.valid) begin
			              n_lkup_reqpkt.lookup=1'b1;
			              n_lkup_reqpkt.hppa=cpu_wr_reqpkt.hppa;	 
			              n_state=WR_LOOKUP_ALLOCATE;
		  	       end
			       else if (cpu_rd_reqpkt.valid) begin 
			              n_lkup_reqpkt.lookup=1'b1;
			              n_lkup_reqpkt.hppa=cpu_rd_reqpkt.hppa;	 
			              n_state=RD_LOOKUP_ALLOCATE;
			       end
			end
		end
		RD_LOOKUP_ALLOCATE: begin
				if(allow_cpu_access) begin 
				      n_allow_cpu_rd_access<=1'b1;
				      n_state<=CHK_WR_ACTIVE;
				end
				else if (tbl_update) begin
				      n_state=RD_TBL_UPDATE;
				end
				//handle inflation later
				//else if (infl)
		end
		WR_LOOKUP_ALLOCATE: begin
				if(allow_cpu_access) begin 
				     n_allow_cpu_wr_access<=1'b1;
				     n_state<=CHK_RD_ACTIVE;
				end
				else if (tbl_update) begin
				     n_state=WR_TBL_UPDATE;
				end
				//handle inflation later
				//else if (infl)
		end
		//The below can be moved to hawk_pgrd_manager, but later it helps
		//to pipeline : look up for pending transactions can be
		//carried out while update table action is pending, move below to other tiny state machine
		//to pipeline 
		RD_TBL_UPDATE:begin
				if(tbl_update_done) begin
					n_allow_cpu_rd_access<=1'b1;
					n_state<=CHK_WR_ACTIVE;
				end
		end
		WR_TBL_UPDATE:begin
				if(tbl_update_done) begin
					n_allow_cpu_wr_access<=1'b1;
					n_state<=CHK_RD_ACTIVE;
				end
		end
	endcase
end

//Flops/State
//state register/output flops
always @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni) begin
		p_state<=IDLE;
		allow_cpu_rd_access<=1'b0;
		allow_cpu_wr_access<=1'b0;
	end
	else begin
		p_state<=n_state;
		allow_cpu_rd_access<=n_allow_cpu_rd_access;
		allow_cpu_wr_access<=n_allow_cpu_wr_access;
	end
end


endmodule
