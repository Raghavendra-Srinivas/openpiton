/////////////////////////////////////////////////////////////////////////////////
//
// Heap Lab Research
// Block : Hawk Page Writer
// 
// Author : Raghavendra Srinivas
// Contact : raghavs@vt.edu	
/////////////////////////////////////////////////////////////////////////////////
// Description: module to handle all page writes from hawk
/////////////////////////////////////////////////////////////////////////////////

module hawk_pg_writer #()
(


);


endmodule
