module hawk_comdecomp (

    
    output wire rdfifo_rdptr_rst, //this would reset read pointer to zero
    input wire  rdfifo_empty,
    input wire  rdfifo_full
);

endmodule
